
module PC ( PC_i, PC_o, clk, rst_n );
  input [31:0] PC_i;
  output [31:0] PC_o;
  input clk, rst_n;
  wire   n1, n2, n3, n4, n5;

  DFFRX1 \PC_o_reg[31]  ( .D(PC_i[31]), .CK(clk), .RN(n5), .Q(PC_o[31]) );
  DFFRX1 \PC_o_reg[29]  ( .D(PC_i[29]), .CK(clk), .RN(n5), .Q(PC_o[29]) );
  DFFRX1 \PC_o_reg[27]  ( .D(PC_i[27]), .CK(clk), .RN(n5), .Q(PC_o[27]) );
  DFFRX1 \PC_o_reg[26]  ( .D(PC_i[26]), .CK(clk), .RN(n5), .Q(PC_o[26]) );
  DFFRX1 \PC_o_reg[25]  ( .D(PC_i[25]), .CK(clk), .RN(n4), .Q(PC_o[25]) );
  DFFRX1 \PC_o_reg[1]  ( .D(PC_i[1]), .CK(clk), .RN(n3), .Q(PC_o[1]) );
  DFFRX1 \PC_o_reg[0]  ( .D(PC_i[0]), .CK(clk), .RN(n3), .Q(PC_o[0]) );
  DFFRX1 \PC_o_reg[24]  ( .D(PC_i[24]), .CK(clk), .RN(n4), .Q(PC_o[24]) );
  DFFRX1 \PC_o_reg[23]  ( .D(PC_i[23]), .CK(clk), .RN(n4), .Q(PC_o[23]) );
  DFFRX1 \PC_o_reg[22]  ( .D(PC_i[22]), .CK(clk), .RN(n4), .Q(PC_o[22]) );
  DFFRX1 \PC_o_reg[21]  ( .D(PC_i[21]), .CK(clk), .RN(n4), .Q(PC_o[21]) );
  DFFRX1 \PC_o_reg[20]  ( .D(PC_i[20]), .CK(clk), .RN(n4), .Q(PC_o[20]) );
  DFFRX1 \PC_o_reg[19]  ( .D(PC_i[19]), .CK(clk), .RN(n4), .Q(PC_o[19]) );
  DFFRX1 \PC_o_reg[18]  ( .D(PC_i[18]), .CK(clk), .RN(n4), .Q(PC_o[18]) );
  DFFRX1 \PC_o_reg[17]  ( .D(PC_i[17]), .CK(clk), .RN(n4), .Q(PC_o[17]) );
  DFFRX1 \PC_o_reg[16]  ( .D(PC_i[16]), .CK(clk), .RN(n4), .Q(PC_o[16]) );
  DFFRX1 \PC_o_reg[15]  ( .D(PC_i[15]), .CK(clk), .RN(n4), .Q(PC_o[15]) );
  DFFRX1 \PC_o_reg[14]  ( .D(PC_i[14]), .CK(clk), .RN(n4), .Q(PC_o[14]) );
  DFFRX1 \PC_o_reg[13]  ( .D(PC_i[13]), .CK(clk), .RN(n4), .Q(PC_o[13]) );
  DFFRX1 \PC_o_reg[12]  ( .D(PC_i[12]), .CK(clk), .RN(n3), .Q(PC_o[12]) );
  DFFRX1 \PC_o_reg[11]  ( .D(PC_i[11]), .CK(clk), .RN(n3), .Q(PC_o[11]) );
  DFFRX1 \PC_o_reg[10]  ( .D(PC_i[10]), .CK(clk), .RN(n3), .Q(PC_o[10]) );
  DFFRX1 \PC_o_reg[9]  ( .D(PC_i[9]), .CK(clk), .RN(n3), .Q(PC_o[9]) );
  DFFRX1 \PC_o_reg[8]  ( .D(PC_i[8]), .CK(clk), .RN(n3), .Q(PC_o[8]) );
  DFFRX1 \PC_o_reg[7]  ( .D(PC_i[7]), .CK(clk), .RN(n3), .Q(PC_o[7]) );
  DFFRX1 \PC_o_reg[6]  ( .D(PC_i[6]), .CK(clk), .RN(n3), .Q(PC_o[6]) );
  DFFRX1 \PC_o_reg[5]  ( .D(PC_i[5]), .CK(clk), .RN(n3), .Q(PC_o[5]) );
  DFFRX1 \PC_o_reg[4]  ( .D(PC_i[4]), .CK(clk), .RN(n3), .Q(PC_o[4]) );
  DFFRX1 \PC_o_reg[3]  ( .D(PC_i[3]), .CK(clk), .RN(n3), .Q(PC_o[3]) );
  DFFRX1 \PC_o_reg[2]  ( .D(PC_i[2]), .CK(clk), .RN(n3), .Q(PC_o[2]) );
  DFFRX1 \PC_o_reg[30]  ( .D(PC_i[30]), .CK(clk), .RN(n5), .Q(PC_o[30]) );
  DFFRX1 \PC_o_reg[28]  ( .D(PC_i[28]), .CK(clk), .RN(n5), .Q(PC_o[28]) );
  CLKBUFX3 U3 ( .A(n1), .Y(n3) );
  CLKBUFX3 U4 ( .A(n1), .Y(n4) );
  CLKBUFX3 U5 ( .A(rst_n), .Y(n1) );
  CLKBUFX3 U6 ( .A(n2), .Y(n5) );
  CLKBUFX3 U7 ( .A(rst_n), .Y(n2) );
endmodule


module Control ( opcode_i, func_i, RegDst_o, Jump_o, Branch_o, MemRead_o, 
        MemToReg_o, ALUOp_o, MemWrite_o, ALUSrc_o, RegWrite_o, jal_o, jr_o );
  input [5:0] opcode_i;
  input [5:0] func_i;
  output [1:0] ALUOp_o;
  output RegDst_o, Jump_o, Branch_o, MemRead_o, MemToReg_o, MemWrite_o,
         ALUSrc_o, RegWrite_o, jal_o, jr_o;
  wire   n6, n7, n8, n9, n10, n11, n12, n4, n5, n13;

  CLKINVX1 U1 ( .A(RegDst_o), .Y(n4) );
  NOR3X1 U2 ( .A(n13), .B(n10), .C(n5), .Y(n8) );
  NAND3BX1 U3 ( .AN(jal_o), .B(n4), .C(n7), .Y(RegWrite_o) );
  CLKINVX1 U4 ( .A(n9), .Y(MemWrite_o) );
  NAND2X1 U5 ( .A(n9), .B(n7), .Y(ALUSrc_o) );
  NOR4X1 U6 ( .A(n10), .B(opcode_i[0]), .C(opcode_i[1]), .D(opcode_i[5]), .Y(
        RegDst_o) );
  NAND3X1 U7 ( .A(n13), .B(n5), .C(opcode_i[2]), .Y(n12) );
  NOR2BX1 U8 ( .AN(n8), .B(opcode_i[5]), .Y(jal_o) );
  NAND4X1 U9 ( .A(opcode_i[5]), .B(opcode_i[1]), .C(opcode_i[3]), .D(n11), .Y(
        n9) );
  NOR3X1 U10 ( .A(n13), .B(opcode_i[4]), .C(opcode_i[2]), .Y(n11) );
  OR3X2 U11 ( .A(opcode_i[3]), .B(opcode_i[4]), .C(opcode_i[2]), .Y(n10) );
  CLKINVX1 U12 ( .A(opcode_i[0]), .Y(n13) );
  CLKINVX1 U13 ( .A(opcode_i[1]), .Y(n5) );
  NAND2X1 U14 ( .A(opcode_i[5]), .B(n8), .Y(n7) );
  NOR4BX1 U15 ( .AN(func_i[3]), .B(n6), .C(func_i[0]), .D(n4), .Y(jr_o) );
  OR4X1 U16 ( .A(func_i[2]), .B(func_i[1]), .C(func_i[5]), .D(func_i[4]), .Y(
        n6) );
  NOR3X1 U17 ( .A(n5), .B(opcode_i[5]), .C(n10), .Y(Jump_o) );
  CLKBUFX3 U18 ( .A(RegDst_o), .Y(ALUOp_o[1]) );
  CLKBUFX3 U19 ( .A(Branch_o), .Y(ALUOp_o[0]) );
  NOR4X1 U20 ( .A(n12), .B(opcode_i[3]), .C(opcode_i[5]), .D(opcode_i[4]), .Y(
        Branch_o) );
  CLKBUFX3 U21 ( .A(MemRead_o), .Y(MemToReg_o) );
  CLKINVX1 U22 ( .A(n7), .Y(MemRead_o) );
endmodule


module MUX2_5b_0 ( data0_i, data1_i, sel_i, data_o );
  input [4:0] data0_i;
  input [4:0] data1_i;
  output [4:0] data_o;
  input sel_i;
  wire   n1;

  CLKINVX1 U1 ( .A(sel_i), .Y(n1) );
  AO22X1 U2 ( .A0(data1_i[2]), .A1(sel_i), .B0(data0_i[2]), .B1(n1), .Y(
        data_o[2]) );
  AO22X1 U3 ( .A0(data1_i[1]), .A1(sel_i), .B0(data0_i[1]), .B1(n1), .Y(
        data_o[1]) );
  AO22X1 U4 ( .A0(sel_i), .A1(data1_i[4]), .B0(data0_i[4]), .B1(n1), .Y(
        data_o[4]) );
  AO22X1 U5 ( .A0(data1_i[0]), .A1(sel_i), .B0(data0_i[0]), .B1(n1), .Y(
        data_o[0]) );
  AO22X1 U6 ( .A0(data1_i[3]), .A1(sel_i), .B0(data0_i[3]), .B1(n1), .Y(
        data_o[3]) );
endmodule


module MUX2_5b_1 ( data0_i, data1_i, sel_i, data_o );
  input [4:0] data0_i;
  input [4:0] data1_i;
  output [4:0] data_o;
  input sel_i;
  wire   n1;

  CLKINVX1 U1 ( .A(sel_i), .Y(n1) );
  AO22X1 U2 ( .A0(data1_i[2]), .A1(sel_i), .B0(data0_i[2]), .B1(n1), .Y(
        data_o[2]) );
  AO22X1 U3 ( .A0(data1_i[1]), .A1(sel_i), .B0(data0_i[1]), .B1(n1), .Y(
        data_o[1]) );
  AO22X1 U4 ( .A0(sel_i), .A1(data1_i[4]), .B0(data0_i[4]), .B1(n1), .Y(
        data_o[4]) );
  AO22X1 U5 ( .A0(data1_i[0]), .A1(sel_i), .B0(data0_i[0]), .B1(n1), .Y(
        data_o[0]) );
  AO22X1 U6 ( .A0(data1_i[3]), .A1(sel_i), .B0(data0_i[3]), .B1(n1), .Y(
        data_o[3]) );
endmodule


module Register ( Reg_R1_i, Reg_R2_i, Reg_W_i, RegWrite_i, WriteData_i, 
        ReadData1_o, ReadData2_o, clk, rst_n );
  input [4:0] Reg_R1_i;
  input [4:0] Reg_R2_i;
  input [4:0] Reg_W_i;
  input [31:0] WriteData_i;
  output [31:0] ReadData1_o;
  output [31:0] ReadData2_o;
  input RegWrite_i, clk, rst_n;
  wire   N467, N468, N469, N470, N471, N472, N473, N474, N475, N476,
         \register[0][31] , \register[0][30] , \register[0][29] ,
         \register[0][28] , \register[0][27] , \register[0][26] ,
         \register[0][25] , \register[0][24] , \register[0][23] ,
         \register[0][22] , \register[0][21] , \register[0][20] ,
         \register[0][19] , \register[0][18] , \register[0][17] ,
         \register[0][16] , \register[0][15] , \register[0][14] ,
         \register[0][13] , \register[0][12] , \register[0][11] ,
         \register[0][10] , \register[0][9] , \register[0][8] ,
         \register[0][7] , \register[0][6] , \register[0][5] ,
         \register[0][4] , \register[0][3] , \register[0][2] ,
         \register[0][1] , \register[0][0] , \register[1][31] ,
         \register[1][30] , \register[1][29] , \register[1][28] ,
         \register[1][27] , \register[1][26] , \register[1][25] ,
         \register[1][24] , \register[1][23] , \register[1][22] ,
         \register[1][21] , \register[1][20] , \register[1][19] ,
         \register[1][18] , \register[1][17] , \register[1][16] ,
         \register[1][15] , \register[1][14] , \register[1][13] ,
         \register[1][12] , \register[1][11] , \register[1][10] ,
         \register[1][9] , \register[1][8] , \register[1][7] ,
         \register[1][6] , \register[1][5] , \register[1][4] ,
         \register[1][3] , \register[1][2] , \register[1][1] ,
         \register[1][0] , \register[2][31] , \register[2][30] ,
         \register[2][29] , \register[2][28] , \register[2][27] ,
         \register[2][26] , \register[2][25] , \register[2][24] ,
         \register[2][23] , \register[2][22] , \register[2][21] ,
         \register[2][20] , \register[2][19] , \register[2][18] ,
         \register[2][17] , \register[2][16] , \register[2][15] ,
         \register[2][14] , \register[2][13] , \register[2][12] ,
         \register[2][11] , \register[2][10] , \register[2][9] ,
         \register[2][8] , \register[2][7] , \register[2][6] ,
         \register[2][5] , \register[2][4] , \register[2][3] ,
         \register[2][2] , \register[2][1] , \register[2][0] ,
         \register[3][31] , \register[3][30] , \register[3][29] ,
         \register[3][28] , \register[3][27] , \register[3][26] ,
         \register[3][25] , \register[3][24] , \register[3][23] ,
         \register[3][22] , \register[3][21] , \register[3][20] ,
         \register[3][19] , \register[3][18] , \register[3][17] ,
         \register[3][16] , \register[3][15] , \register[3][14] ,
         \register[3][13] , \register[3][12] , \register[3][11] ,
         \register[3][10] , \register[3][9] , \register[3][8] ,
         \register[3][7] , \register[3][6] , \register[3][5] ,
         \register[3][4] , \register[3][3] , \register[3][2] ,
         \register[3][1] , \register[3][0] , \register[4][31] ,
         \register[4][30] , \register[4][29] , \register[4][28] ,
         \register[4][27] , \register[4][26] , \register[4][25] ,
         \register[4][24] , \register[4][23] , \register[4][22] ,
         \register[4][21] , \register[4][20] , \register[4][19] ,
         \register[4][18] , \register[4][17] , \register[4][16] ,
         \register[4][15] , \register[4][14] , \register[4][13] ,
         \register[4][12] , \register[4][11] , \register[4][10] ,
         \register[4][9] , \register[4][8] , \register[4][7] ,
         \register[4][6] , \register[4][5] , \register[4][4] ,
         \register[4][3] , \register[4][2] , \register[4][1] ,
         \register[4][0] , \register[5][31] , \register[5][30] ,
         \register[5][29] , \register[5][28] , \register[5][27] ,
         \register[5][26] , \register[5][25] , \register[5][24] ,
         \register[5][23] , \register[5][22] , \register[5][21] ,
         \register[5][20] , \register[5][19] , \register[5][18] ,
         \register[5][17] , \register[5][16] , \register[5][15] ,
         \register[5][14] , \register[5][13] , \register[5][12] ,
         \register[5][11] , \register[5][10] , \register[5][9] ,
         \register[5][8] , \register[5][7] , \register[5][6] ,
         \register[5][5] , \register[5][4] , \register[5][3] ,
         \register[5][2] , \register[5][1] , \register[5][0] ,
         \register[6][31] , \register[6][30] , \register[6][29] ,
         \register[6][28] , \register[6][27] , \register[6][26] ,
         \register[6][25] , \register[6][24] , \register[6][23] ,
         \register[6][22] , \register[6][21] , \register[6][20] ,
         \register[6][19] , \register[6][18] , \register[6][17] ,
         \register[6][16] , \register[6][15] , \register[6][14] ,
         \register[6][13] , \register[6][12] , \register[6][11] ,
         \register[6][10] , \register[6][9] , \register[6][8] ,
         \register[6][7] , \register[6][6] , \register[6][5] ,
         \register[6][4] , \register[6][3] , \register[6][2] ,
         \register[6][1] , \register[6][0] , \register[7][31] ,
         \register[7][30] , \register[7][29] , \register[7][28] ,
         \register[7][27] , \register[7][26] , \register[7][25] ,
         \register[7][24] , \register[7][23] , \register[7][22] ,
         \register[7][21] , \register[7][20] , \register[7][19] ,
         \register[7][18] , \register[7][17] , \register[7][16] ,
         \register[7][15] , \register[7][14] , \register[7][13] ,
         \register[7][12] , \register[7][11] , \register[7][10] ,
         \register[7][9] , \register[7][8] , \register[7][7] ,
         \register[7][6] , \register[7][5] , \register[7][4] ,
         \register[7][3] , \register[7][2] , \register[7][1] ,
         \register[7][0] , \register[8][31] , \register[8][30] ,
         \register[8][29] , \register[8][28] , \register[8][27] ,
         \register[8][26] , \register[8][25] , \register[8][24] ,
         \register[8][23] , \register[8][22] , \register[8][21] ,
         \register[8][20] , \register[8][19] , \register[8][18] ,
         \register[8][17] , \register[8][16] , \register[8][15] ,
         \register[8][14] , \register[8][13] , \register[8][12] ,
         \register[8][11] , \register[8][10] , \register[8][9] ,
         \register[8][8] , \register[8][7] , \register[8][6] ,
         \register[8][5] , \register[8][4] , \register[8][3] ,
         \register[8][2] , \register[8][1] , \register[8][0] ,
         \register[9][31] , \register[9][30] , \register[9][29] ,
         \register[9][28] , \register[9][27] , \register[9][26] ,
         \register[9][25] , \register[9][24] , \register[9][23] ,
         \register[9][22] , \register[9][21] , \register[9][20] ,
         \register[9][19] , \register[9][18] , \register[9][17] ,
         \register[9][16] , \register[9][15] , \register[9][14] ,
         \register[9][13] , \register[9][12] , \register[9][11] ,
         \register[9][10] , \register[9][9] , \register[9][8] ,
         \register[9][7] , \register[9][6] , \register[9][5] ,
         \register[9][4] , \register[9][3] , \register[9][2] ,
         \register[9][1] , \register[9][0] , \register[10][31] ,
         \register[10][30] , \register[10][29] , \register[10][28] ,
         \register[10][27] , \register[10][26] , \register[10][25] ,
         \register[10][24] , \register[10][23] , \register[10][22] ,
         \register[10][21] , \register[10][20] , \register[10][19] ,
         \register[10][18] , \register[10][17] , \register[10][16] ,
         \register[10][15] , \register[10][14] , \register[10][13] ,
         \register[10][12] , \register[10][11] , \register[10][10] ,
         \register[10][9] , \register[10][8] , \register[10][7] ,
         \register[10][6] , \register[10][5] , \register[10][4] ,
         \register[10][3] , \register[10][2] , \register[10][1] ,
         \register[10][0] , \register[11][31] , \register[11][30] ,
         \register[11][29] , \register[11][28] , \register[11][27] ,
         \register[11][26] , \register[11][25] , \register[11][24] ,
         \register[11][23] , \register[11][22] , \register[11][21] ,
         \register[11][20] , \register[11][19] , \register[11][18] ,
         \register[11][17] , \register[11][16] , \register[11][15] ,
         \register[11][14] , \register[11][13] , \register[11][12] ,
         \register[11][11] , \register[11][10] , \register[11][9] ,
         \register[11][8] , \register[11][7] , \register[11][6] ,
         \register[11][5] , \register[11][4] , \register[11][3] ,
         \register[11][2] , \register[11][1] , \register[11][0] ,
         \register[12][31] , \register[12][30] , \register[12][29] ,
         \register[12][28] , \register[12][27] , \register[12][26] ,
         \register[12][25] , \register[12][24] , \register[12][23] ,
         \register[12][22] , \register[12][21] , \register[12][20] ,
         \register[12][19] , \register[12][18] , \register[12][17] ,
         \register[12][16] , \register[12][15] , \register[12][14] ,
         \register[12][13] , \register[12][12] , \register[12][11] ,
         \register[12][10] , \register[12][9] , \register[12][8] ,
         \register[12][7] , \register[12][6] , \register[12][5] ,
         \register[12][4] , \register[12][3] , \register[12][2] ,
         \register[12][1] , \register[12][0] , \register[13][31] ,
         \register[13][30] , \register[13][29] , \register[13][28] ,
         \register[13][27] , \register[13][26] , \register[13][25] ,
         \register[13][24] , \register[13][23] , \register[13][22] ,
         \register[13][21] , \register[13][20] , \register[13][19] ,
         \register[13][18] , \register[13][17] , \register[13][16] ,
         \register[13][15] , \register[13][14] , \register[13][13] ,
         \register[13][12] , \register[13][11] , \register[13][10] ,
         \register[13][9] , \register[13][8] , \register[13][7] ,
         \register[13][6] , \register[13][5] , \register[13][4] ,
         \register[13][3] , \register[13][2] , \register[13][1] ,
         \register[13][0] , \register[14][31] , \register[14][30] ,
         \register[14][29] , \register[14][28] , \register[14][27] ,
         \register[14][26] , \register[14][25] , \register[14][24] ,
         \register[14][23] , \register[14][22] , \register[14][21] ,
         \register[14][20] , \register[14][19] , \register[14][18] ,
         \register[14][17] , \register[14][16] , \register[14][15] ,
         \register[14][14] , \register[14][13] , \register[14][12] ,
         \register[14][11] , \register[14][10] , \register[14][9] ,
         \register[14][8] , \register[14][7] , \register[14][6] ,
         \register[14][5] , \register[14][4] , \register[14][3] ,
         \register[14][2] , \register[14][1] , \register[14][0] ,
         \register[15][31] , \register[15][30] , \register[15][29] ,
         \register[15][28] , \register[15][27] , \register[15][26] ,
         \register[15][25] , \register[15][24] , \register[15][23] ,
         \register[15][22] , \register[15][21] , \register[15][20] ,
         \register[15][19] , \register[15][18] , \register[15][17] ,
         \register[15][16] , \register[15][15] , \register[15][14] ,
         \register[15][13] , \register[15][12] , \register[15][11] ,
         \register[15][10] , \register[15][9] , \register[15][8] ,
         \register[15][7] , \register[15][6] , \register[15][5] ,
         \register[15][4] , \register[15][3] , \register[15][2] ,
         \register[15][1] , \register[15][0] , \register[16][31] ,
         \register[16][30] , \register[16][29] , \register[16][28] ,
         \register[16][27] , \register[16][26] , \register[16][25] ,
         \register[16][24] , \register[16][23] , \register[16][22] ,
         \register[16][21] , \register[16][20] , \register[16][19] ,
         \register[16][18] , \register[16][17] , \register[16][16] ,
         \register[16][15] , \register[16][14] , \register[16][13] ,
         \register[16][12] , \register[16][11] , \register[16][10] ,
         \register[16][9] , \register[16][8] , \register[16][7] ,
         \register[16][6] , \register[16][5] , \register[16][4] ,
         \register[16][3] , \register[16][2] , \register[16][1] ,
         \register[16][0] , \register[17][31] , \register[17][30] ,
         \register[17][29] , \register[17][28] , \register[17][27] ,
         \register[17][26] , \register[17][25] , \register[17][24] ,
         \register[17][23] , \register[17][22] , \register[17][21] ,
         \register[17][20] , \register[17][19] , \register[17][18] ,
         \register[17][17] , \register[17][16] , \register[17][15] ,
         \register[17][14] , \register[17][13] , \register[17][12] ,
         \register[17][11] , \register[17][10] , \register[17][9] ,
         \register[17][8] , \register[17][7] , \register[17][6] ,
         \register[17][5] , \register[17][4] , \register[17][3] ,
         \register[17][2] , \register[17][1] , \register[17][0] ,
         \register[18][31] , \register[18][30] , \register[18][29] ,
         \register[18][28] , \register[18][27] , \register[18][26] ,
         \register[18][25] , \register[18][24] , \register[18][23] ,
         \register[18][22] , \register[18][21] , \register[18][20] ,
         \register[18][19] , \register[18][18] , \register[18][17] ,
         \register[18][16] , \register[18][15] , \register[18][14] ,
         \register[18][13] , \register[18][12] , \register[18][11] ,
         \register[18][10] , \register[18][9] , \register[18][8] ,
         \register[18][7] , \register[18][6] , \register[18][5] ,
         \register[18][4] , \register[18][3] , \register[18][2] ,
         \register[18][1] , \register[18][0] , \register[19][31] ,
         \register[19][30] , \register[19][29] , \register[19][28] ,
         \register[19][27] , \register[19][26] , \register[19][25] ,
         \register[19][24] , \register[19][23] , \register[19][22] ,
         \register[19][21] , \register[19][20] , \register[19][19] ,
         \register[19][18] , \register[19][17] , \register[19][16] ,
         \register[19][15] , \register[19][14] , \register[19][13] ,
         \register[19][12] , \register[19][11] , \register[19][10] ,
         \register[19][9] , \register[19][8] , \register[19][7] ,
         \register[19][6] , \register[19][5] , \register[19][4] ,
         \register[19][3] , \register[19][2] , \register[19][1] ,
         \register[19][0] , \register[20][31] , \register[20][30] ,
         \register[20][29] , \register[20][28] , \register[20][27] ,
         \register[20][26] , \register[20][25] , \register[20][24] ,
         \register[20][23] , \register[20][22] , \register[20][21] ,
         \register[20][20] , \register[20][19] , \register[20][18] ,
         \register[20][17] , \register[20][16] , \register[20][15] ,
         \register[20][14] , \register[20][13] , \register[20][12] ,
         \register[20][11] , \register[20][10] , \register[20][9] ,
         \register[20][8] , \register[20][7] , \register[20][6] ,
         \register[20][5] , \register[20][4] , \register[20][3] ,
         \register[20][2] , \register[20][1] , \register[20][0] ,
         \register[21][31] , \register[21][30] , \register[21][29] ,
         \register[21][28] , \register[21][27] , \register[21][26] ,
         \register[21][25] , \register[21][24] , \register[21][23] ,
         \register[21][22] , \register[21][21] , \register[21][20] ,
         \register[21][19] , \register[21][18] , \register[21][17] ,
         \register[21][16] , \register[21][15] , \register[21][14] ,
         \register[21][13] , \register[21][12] , \register[21][11] ,
         \register[21][10] , \register[21][9] , \register[21][8] ,
         \register[21][7] , \register[21][6] , \register[21][5] ,
         \register[21][4] , \register[21][3] , \register[21][2] ,
         \register[21][1] , \register[21][0] , \register[22][31] ,
         \register[22][30] , \register[22][29] , \register[22][28] ,
         \register[22][27] , \register[22][26] , \register[22][25] ,
         \register[22][24] , \register[22][23] , \register[22][22] ,
         \register[22][21] , \register[22][20] , \register[22][19] ,
         \register[22][18] , \register[22][17] , \register[22][16] ,
         \register[22][15] , \register[22][14] , \register[22][13] ,
         \register[22][12] , \register[22][11] , \register[22][10] ,
         \register[22][9] , \register[22][8] , \register[22][7] ,
         \register[22][6] , \register[22][5] , \register[22][4] ,
         \register[22][3] , \register[22][2] , \register[22][1] ,
         \register[22][0] , \register[23][31] , \register[23][30] ,
         \register[23][29] , \register[23][28] , \register[23][27] ,
         \register[23][26] , \register[23][25] , \register[23][24] ,
         \register[23][23] , \register[23][22] , \register[23][21] ,
         \register[23][20] , \register[23][19] , \register[23][18] ,
         \register[23][17] , \register[23][16] , \register[23][15] ,
         \register[23][14] , \register[23][13] , \register[23][12] ,
         \register[23][11] , \register[23][10] , \register[23][9] ,
         \register[23][8] , \register[23][7] , \register[23][6] ,
         \register[23][5] , \register[23][4] , \register[23][3] ,
         \register[23][2] , \register[23][1] , \register[23][0] ,
         \register[24][31] , \register[24][30] , \register[24][29] ,
         \register[24][28] , \register[24][27] , \register[24][26] ,
         \register[24][25] , \register[24][24] , \register[24][23] ,
         \register[24][22] , \register[24][21] , \register[24][20] ,
         \register[24][19] , \register[24][18] , \register[24][17] ,
         \register[24][16] , \register[24][15] , \register[24][14] ,
         \register[24][13] , \register[24][12] , \register[24][11] ,
         \register[24][10] , \register[24][9] , \register[24][8] ,
         \register[24][7] , \register[24][6] , \register[24][5] ,
         \register[24][4] , \register[24][3] , \register[24][2] ,
         \register[24][1] , \register[24][0] , \register[25][31] ,
         \register[25][30] , \register[25][29] , \register[25][28] ,
         \register[25][27] , \register[25][26] , \register[25][25] ,
         \register[25][24] , \register[25][23] , \register[25][22] ,
         \register[25][21] , \register[25][20] , \register[25][19] ,
         \register[25][18] , \register[25][17] , \register[25][16] ,
         \register[25][15] , \register[25][14] , \register[25][13] ,
         \register[25][12] , \register[25][11] , \register[25][10] ,
         \register[25][9] , \register[25][8] , \register[25][7] ,
         \register[25][6] , \register[25][5] , \register[25][4] ,
         \register[25][3] , \register[25][2] , \register[25][1] ,
         \register[25][0] , \register[26][31] , \register[26][30] ,
         \register[26][29] , \register[26][28] , \register[26][27] ,
         \register[26][26] , \register[26][25] , \register[26][24] ,
         \register[26][23] , \register[26][22] , \register[26][21] ,
         \register[26][20] , \register[26][19] , \register[26][18] ,
         \register[26][17] , \register[26][16] , \register[26][15] ,
         \register[26][14] , \register[26][13] , \register[26][12] ,
         \register[26][11] , \register[26][10] , \register[26][9] ,
         \register[26][8] , \register[26][7] , \register[26][6] ,
         \register[26][5] , \register[26][4] , \register[26][3] ,
         \register[26][2] , \register[26][1] , \register[26][0] ,
         \register[27][31] , \register[27][30] , \register[27][29] ,
         \register[27][28] , \register[27][27] , \register[27][26] ,
         \register[27][25] , \register[27][24] , \register[27][23] ,
         \register[27][22] , \register[27][21] , \register[27][20] ,
         \register[27][19] , \register[27][18] , \register[27][17] ,
         \register[27][16] , \register[27][15] , \register[27][14] ,
         \register[27][13] , \register[27][12] , \register[27][11] ,
         \register[27][10] , \register[27][9] , \register[27][8] ,
         \register[27][7] , \register[27][6] , \register[27][5] ,
         \register[27][4] , \register[27][3] , \register[27][2] ,
         \register[27][1] , \register[27][0] , \register[28][31] ,
         \register[28][30] , \register[28][29] , \register[28][28] ,
         \register[28][27] , \register[28][26] , \register[28][25] ,
         \register[28][24] , \register[28][23] , \register[28][22] ,
         \register[28][21] , \register[28][20] , \register[28][19] ,
         \register[28][18] , \register[28][17] , \register[28][16] ,
         \register[28][15] , \register[28][14] , \register[28][13] ,
         \register[28][12] , \register[28][11] , \register[28][10] ,
         \register[28][9] , \register[28][8] , \register[28][7] ,
         \register[28][6] , \register[28][5] , \register[28][4] ,
         \register[28][3] , \register[28][2] , \register[28][1] ,
         \register[28][0] , \register[29][31] , \register[29][30] ,
         \register[29][29] , \register[29][28] , \register[29][27] ,
         \register[29][26] , \register[29][25] , \register[29][24] ,
         \register[29][23] , \register[29][22] , \register[29][21] ,
         \register[29][20] , \register[29][19] , \register[29][18] ,
         \register[29][17] , \register[29][16] , \register[29][15] ,
         \register[29][14] , \register[29][13] , \register[29][12] ,
         \register[29][11] , \register[29][10] , \register[29][9] ,
         \register[29][8] , \register[29][7] , \register[29][6] ,
         \register[29][5] , \register[29][4] , \register[29][3] ,
         \register[29][2] , \register[29][1] , \register[29][0] ,
         \register[30][31] , \register[30][30] , \register[30][29] ,
         \register[30][28] , \register[30][27] , \register[30][26] ,
         \register[30][25] , \register[30][24] , \register[30][23] ,
         \register[30][22] , \register[30][21] , \register[30][20] ,
         \register[30][19] , \register[30][18] , \register[30][17] ,
         \register[30][16] , \register[30][15] , \register[30][14] ,
         \register[30][13] , \register[30][12] , \register[30][11] ,
         \register[30][10] , \register[30][9] , \register[30][8] ,
         \register[30][7] , \register[30][6] , \register[30][5] ,
         \register[30][4] , \register[30][3] , \register[30][2] ,
         \register[30][1] , \register[30][0] , \register[31][31] ,
         \register[31][30] , \register[31][29] , \register[31][28] ,
         \register[31][27] , \register[31][26] , \register[31][25] ,
         \register[31][24] , \register[31][23] , \register[31][22] ,
         \register[31][21] , \register[31][20] , \register[31][19] ,
         \register[31][18] , \register[31][17] , \register[31][16] ,
         \register[31][15] , \register[31][14] , \register[31][13] ,
         \register[31][12] , \register[31][11] , \register[31][10] ,
         \register[31][9] , \register[31][8] , \register[31][7] ,
         \register[31][6] , \register[31][5] , \register[31][4] ,
         \register[31][3] , \register[31][2] , \register[31][1] ,
         \register[31][0] , n69, n70, n104, n138, n172, n206, n240, n274, n308,
         n342, n607, n872, n873, n907, n941, n975, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355;
  assign N467 = Reg_R1_i[0];
  assign N468 = Reg_R1_i[1];
  assign N469 = Reg_R1_i[2];
  assign N470 = Reg_R1_i[3];
  assign N471 = Reg_R1_i[4];
  assign N472 = Reg_R2_i[0];
  assign N473 = Reg_R2_i[1];
  assign N474 = Reg_R2_i[2];
  assign N475 = Reg_R2_i[3];
  assign N476 = Reg_R2_i[4];

  DFFRX1 \register_reg[3][31]  ( .D(n1140), .CK(clk), .RN(n2280), .Q(
        \register[3][31] ) );
  DFFRX1 \register_reg[3][30]  ( .D(n1141), .CK(clk), .RN(n2280), .Q(
        \register[3][30] ) );
  DFFRX1 \register_reg[3][29]  ( .D(n1142), .CK(clk), .RN(n2280), .Q(
        \register[3][29] ) );
  DFFRX1 \register_reg[3][28]  ( .D(n1143), .CK(clk), .RN(n2280), .Q(
        \register[3][28] ) );
  DFFRX1 \register_reg[3][27]  ( .D(n1144), .CK(clk), .RN(n2280), .Q(
        \register[3][27] ) );
  DFFRX1 \register_reg[3][26]  ( .D(n1145), .CK(clk), .RN(n2279), .Q(
        \register[3][26] ) );
  DFFRX1 \register_reg[3][25]  ( .D(n1146), .CK(clk), .RN(n2279), .Q(
        \register[3][25] ) );
  DFFRX1 \register_reg[3][24]  ( .D(n1147), .CK(clk), .RN(n2279), .Q(
        \register[3][24] ) );
  DFFRX1 \register_reg[3][23]  ( .D(n1148), .CK(clk), .RN(n2279), .Q(
        \register[3][23] ) );
  DFFRX1 \register_reg[3][22]  ( .D(n1149), .CK(clk), .RN(n2279), .Q(
        \register[3][22] ) );
  DFFRX1 \register_reg[3][21]  ( .D(n1150), .CK(clk), .RN(n2279), .Q(
        \register[3][21] ) );
  DFFRX1 \register_reg[3][20]  ( .D(n1151), .CK(clk), .RN(n2279), .Q(
        \register[3][20] ) );
  DFFRX1 \register_reg[3][19]  ( .D(n1152), .CK(clk), .RN(n2279), .Q(
        \register[3][19] ) );
  DFFRX1 \register_reg[3][18]  ( .D(n1153), .CK(clk), .RN(n2279), .Q(
        \register[3][18] ) );
  DFFRX1 \register_reg[3][17]  ( .D(n1154), .CK(clk), .RN(n2279), .Q(
        \register[3][17] ) );
  DFFRX1 \register_reg[3][16]  ( .D(n1155), .CK(clk), .RN(n2279), .Q(
        \register[3][16] ) );
  DFFRX1 \register_reg[3][15]  ( .D(n1156), .CK(clk), .RN(n2279), .Q(
        \register[3][15] ) );
  DFFRX1 \register_reg[3][14]  ( .D(n1157), .CK(clk), .RN(n2279), .Q(
        \register[3][14] ) );
  DFFRX1 \register_reg[3][13]  ( .D(n1158), .CK(clk), .RN(n2278), .Q(
        \register[3][13] ) );
  DFFRX1 \register_reg[3][12]  ( .D(n1159), .CK(clk), .RN(n2278), .Q(
        \register[3][12] ) );
  DFFRX1 \register_reg[3][11]  ( .D(n1160), .CK(clk), .RN(n2278), .Q(
        \register[3][11] ) );
  DFFRX1 \register_reg[3][10]  ( .D(n1161), .CK(clk), .RN(n2278), .Q(
        \register[3][10] ) );
  DFFRX1 \register_reg[3][9]  ( .D(n1162), .CK(clk), .RN(n2278), .Q(
        \register[3][9] ) );
  DFFRX1 \register_reg[7][31]  ( .D(n1268), .CK(clk), .RN(n2270), .Q(
        \register[7][31] ) );
  DFFRX1 \register_reg[7][30]  ( .D(n1269), .CK(clk), .RN(n2270), .Q(
        \register[7][30] ) );
  DFFRX1 \register_reg[7][29]  ( .D(n1270), .CK(clk), .RN(n2270), .Q(
        \register[7][29] ) );
  DFFRX1 \register_reg[7][28]  ( .D(n1271), .CK(clk), .RN(n2270), .Q(
        \register[7][28] ) );
  DFFRX1 \register_reg[7][27]  ( .D(n1272), .CK(clk), .RN(n2270), .Q(
        \register[7][27] ) );
  DFFRX1 \register_reg[7][26]  ( .D(n1273), .CK(clk), .RN(n2270), .Q(
        \register[7][26] ) );
  DFFRX1 \register_reg[7][25]  ( .D(n1274), .CK(clk), .RN(n2270), .Q(
        \register[7][25] ) );
  DFFRX1 \register_reg[7][24]  ( .D(n1275), .CK(clk), .RN(n2269), .Q(
        \register[7][24] ) );
  DFFRX1 \register_reg[7][23]  ( .D(n1276), .CK(clk), .RN(n2269), .Q(
        \register[7][23] ) );
  DFFRX1 \register_reg[7][22]  ( .D(n1277), .CK(clk), .RN(n2269), .Q(
        \register[7][22] ) );
  DFFRX1 \register_reg[7][21]  ( .D(n1278), .CK(clk), .RN(n2269), .Q(
        \register[7][21] ) );
  DFFRX1 \register_reg[7][20]  ( .D(n1279), .CK(clk), .RN(n2269), .Q(
        \register[7][20] ) );
  DFFRX1 \register_reg[7][19]  ( .D(n1280), .CK(clk), .RN(n2269), .Q(
        \register[7][19] ) );
  DFFRX1 \register_reg[7][18]  ( .D(n1281), .CK(clk), .RN(n2269), .Q(
        \register[7][18] ) );
  DFFRX1 \register_reg[7][17]  ( .D(n1282), .CK(clk), .RN(n2269), .Q(
        \register[7][17] ) );
  DFFRX1 \register_reg[7][16]  ( .D(n1283), .CK(clk), .RN(n2269), .Q(
        \register[7][16] ) );
  DFFRX1 \register_reg[7][15]  ( .D(n1284), .CK(clk), .RN(n2269), .Q(
        \register[7][15] ) );
  DFFRX1 \register_reg[7][14]  ( .D(n1285), .CK(clk), .RN(n2269), .Q(
        \register[7][14] ) );
  DFFRX1 \register_reg[7][13]  ( .D(n1286), .CK(clk), .RN(n2269), .Q(
        \register[7][13] ) );
  DFFRX1 \register_reg[7][12]  ( .D(n1287), .CK(clk), .RN(n2269), .Q(
        \register[7][12] ) );
  DFFRX1 \register_reg[7][11]  ( .D(n1288), .CK(clk), .RN(n2268), .Q(
        \register[7][11] ) );
  DFFRX1 \register_reg[7][10]  ( .D(n1289), .CK(clk), .RN(n2268), .Q(
        \register[7][10] ) );
  DFFRX1 \register_reg[7][9]  ( .D(n1290), .CK(clk), .RN(n2268), .Q(
        \register[7][9] ) );
  DFFRX1 \register_reg[11][31]  ( .D(n1396), .CK(clk), .RN(n2260), .Q(
        \register[11][31] ) );
  DFFRX1 \register_reg[11][30]  ( .D(n1397), .CK(clk), .RN(n2260), .Q(
        \register[11][30] ) );
  DFFRX1 \register_reg[11][29]  ( .D(n1398), .CK(clk), .RN(n2260), .Q(
        \register[11][29] ) );
  DFFRX1 \register_reg[11][28]  ( .D(n1399), .CK(clk), .RN(n2260), .Q(
        \register[11][28] ) );
  DFFRX1 \register_reg[11][27]  ( .D(n1400), .CK(clk), .RN(n2260), .Q(
        \register[11][27] ) );
  DFFRX1 \register_reg[11][26]  ( .D(n1401), .CK(clk), .RN(n2260), .Q(
        \register[11][26] ) );
  DFFRX1 \register_reg[11][25]  ( .D(n1402), .CK(clk), .RN(n2260), .Q(
        \register[11][25] ) );
  DFFRX1 \register_reg[11][24]  ( .D(n1403), .CK(clk), .RN(n2260), .Q(
        \register[11][24] ) );
  DFFRX1 \register_reg[11][23]  ( .D(n1404), .CK(clk), .RN(n2260), .Q(
        \register[11][23] ) );
  DFFRX1 \register_reg[11][22]  ( .D(n1405), .CK(clk), .RN(n2259), .Q(
        \register[11][22] ) );
  DFFRX1 \register_reg[11][21]  ( .D(n1406), .CK(clk), .RN(n2259), .Q(
        \register[11][21] ) );
  DFFRX1 \register_reg[11][20]  ( .D(n1407), .CK(clk), .RN(n2259), .Q(
        \register[11][20] ) );
  DFFRX1 \register_reg[11][19]  ( .D(n1408), .CK(clk), .RN(n2259), .Q(
        \register[11][19] ) );
  DFFRX1 \register_reg[11][18]  ( .D(n1409), .CK(clk), .RN(n2259), .Q(
        \register[11][18] ) );
  DFFRX1 \register_reg[11][17]  ( .D(n1410), .CK(clk), .RN(n2259), .Q(
        \register[11][17] ) );
  DFFRX1 \register_reg[11][16]  ( .D(n1411), .CK(clk), .RN(n2259), .Q(
        \register[11][16] ) );
  DFFRX1 \register_reg[11][15]  ( .D(n1412), .CK(clk), .RN(n2259), .Q(
        \register[11][15] ) );
  DFFRX1 \register_reg[11][14]  ( .D(n1413), .CK(clk), .RN(n2259), .Q(
        \register[11][14] ) );
  DFFRX1 \register_reg[11][13]  ( .D(n1414), .CK(clk), .RN(n2259), .Q(
        \register[11][13] ) );
  DFFRX1 \register_reg[11][12]  ( .D(n1415), .CK(clk), .RN(n2259), .Q(
        \register[11][12] ) );
  DFFRX1 \register_reg[11][11]  ( .D(n1416), .CK(clk), .RN(n2259), .Q(
        \register[11][11] ) );
  DFFRX1 \register_reg[11][10]  ( .D(n1417), .CK(clk), .RN(n2259), .Q(
        \register[11][10] ) );
  DFFRX1 \register_reg[11][9]  ( .D(n1418), .CK(clk), .RN(n2258), .Q(
        \register[11][9] ) );
  DFFRX1 \register_reg[15][31]  ( .D(n1524), .CK(clk), .RN(n2250), .Q(
        \register[15][31] ) );
  DFFRX1 \register_reg[15][30]  ( .D(n1525), .CK(clk), .RN(n2250), .Q(
        \register[15][30] ) );
  DFFRX1 \register_reg[15][29]  ( .D(n1526), .CK(clk), .RN(n2250), .Q(
        \register[15][29] ) );
  DFFRX1 \register_reg[15][28]  ( .D(n1527), .CK(clk), .RN(n2250), .Q(
        \register[15][28] ) );
  DFFRX1 \register_reg[15][27]  ( .D(n1528), .CK(clk), .RN(n2250), .Q(
        \register[15][27] ) );
  DFFRX1 \register_reg[15][26]  ( .D(n1529), .CK(clk), .RN(n2250), .Q(
        \register[15][26] ) );
  DFFRX1 \register_reg[15][25]  ( .D(n1530), .CK(clk), .RN(n2250), .Q(
        \register[15][25] ) );
  DFFRX1 \register_reg[15][24]  ( .D(n1531), .CK(clk), .RN(n2250), .Q(
        \register[15][24] ) );
  DFFRX1 \register_reg[15][23]  ( .D(n1532), .CK(clk), .RN(n2250), .Q(
        \register[15][23] ) );
  DFFRX1 \register_reg[15][22]  ( .D(n1533), .CK(clk), .RN(n2250), .Q(
        \register[15][22] ) );
  DFFRX1 \register_reg[15][21]  ( .D(n1534), .CK(clk), .RN(n2250), .Q(
        \register[15][21] ) );
  DFFRX1 \register_reg[15][20]  ( .D(n1535), .CK(clk), .RN(n2249), .Q(
        \register[15][20] ) );
  DFFRX1 \register_reg[15][19]  ( .D(n1536), .CK(clk), .RN(n2249), .Q(
        \register[15][19] ) );
  DFFRX1 \register_reg[15][18]  ( .D(n1537), .CK(clk), .RN(n2249), .Q(
        \register[15][18] ) );
  DFFRX1 \register_reg[15][17]  ( .D(n1538), .CK(clk), .RN(n2249), .Q(
        \register[15][17] ) );
  DFFRX1 \register_reg[15][16]  ( .D(n1539), .CK(clk), .RN(n2249), .Q(
        \register[15][16] ) );
  DFFRX1 \register_reg[15][15]  ( .D(n1540), .CK(clk), .RN(n2249), .Q(
        \register[15][15] ) );
  DFFRX1 \register_reg[15][14]  ( .D(n1541), .CK(clk), .RN(n2249), .Q(
        \register[15][14] ) );
  DFFRX1 \register_reg[15][13]  ( .D(n1542), .CK(clk), .RN(n2249), .Q(
        \register[15][13] ) );
  DFFRX1 \register_reg[15][12]  ( .D(n1543), .CK(clk), .RN(n2249), .Q(
        \register[15][12] ) );
  DFFRX1 \register_reg[15][11]  ( .D(n1544), .CK(clk), .RN(n2249), .Q(
        \register[15][11] ) );
  DFFRX1 \register_reg[15][10]  ( .D(n1545), .CK(clk), .RN(n2249), .Q(
        \register[15][10] ) );
  DFFRX1 \register_reg[15][9]  ( .D(n1546), .CK(clk), .RN(n2249), .Q(
        \register[15][9] ) );
  DFFRX1 \register_reg[19][31]  ( .D(n1652), .CK(clk), .RN(n2240), .Q(
        \register[19][31] ) );
  DFFRX1 \register_reg[19][30]  ( .D(n1653), .CK(clk), .RN(n2240), .Q(
        \register[19][30] ) );
  DFFRX1 \register_reg[19][29]  ( .D(n1654), .CK(clk), .RN(n2240), .Q(
        \register[19][29] ) );
  DFFRX1 \register_reg[19][28]  ( .D(n1655), .CK(clk), .RN(n2240), .Q(
        \register[19][28] ) );
  DFFRX1 \register_reg[19][27]  ( .D(n1656), .CK(clk), .RN(n2240), .Q(
        \register[19][27] ) );
  DFFRX1 \register_reg[19][26]  ( .D(n1657), .CK(clk), .RN(n2240), .Q(
        \register[19][26] ) );
  DFFRX1 \register_reg[19][25]  ( .D(n1658), .CK(clk), .RN(n2240), .Q(
        \register[19][25] ) );
  DFFRX1 \register_reg[19][24]  ( .D(n1659), .CK(clk), .RN(n2240), .Q(
        \register[19][24] ) );
  DFFRX1 \register_reg[19][23]  ( .D(n1660), .CK(clk), .RN(n2240), .Q(
        \register[19][23] ) );
  DFFRX1 \register_reg[19][22]  ( .D(n1661), .CK(clk), .RN(n2240), .Q(
        \register[19][22] ) );
  DFFRX1 \register_reg[19][21]  ( .D(n1662), .CK(clk), .RN(n2240), .Q(
        \register[19][21] ) );
  DFFRX1 \register_reg[19][20]  ( .D(n1663), .CK(clk), .RN(n2240), .Q(
        \register[19][20] ) );
  DFFRX1 \register_reg[19][19]  ( .D(n1664), .CK(clk), .RN(n2240), .Q(
        \register[19][19] ) );
  DFFRX1 \register_reg[19][18]  ( .D(n1665), .CK(clk), .RN(n2239), .Q(
        \register[19][18] ) );
  DFFRX1 \register_reg[19][17]  ( .D(n1666), .CK(clk), .RN(n2239), .Q(
        \register[19][17] ) );
  DFFRX1 \register_reg[19][16]  ( .D(n1667), .CK(clk), .RN(n2239), .Q(
        \register[19][16] ) );
  DFFRX1 \register_reg[19][15]  ( .D(n1668), .CK(clk), .RN(n2239), .Q(
        \register[19][15] ) );
  DFFRX1 \register_reg[19][14]  ( .D(n1669), .CK(clk), .RN(n2239), .Q(
        \register[19][14] ) );
  DFFRX1 \register_reg[19][13]  ( .D(n1670), .CK(clk), .RN(n2239), .Q(
        \register[19][13] ) );
  DFFRX1 \register_reg[19][12]  ( .D(n1671), .CK(clk), .RN(n2239), .Q(
        \register[19][12] ) );
  DFFRX1 \register_reg[19][11]  ( .D(n1672), .CK(clk), .RN(n2239), .Q(
        \register[19][11] ) );
  DFFRX1 \register_reg[19][10]  ( .D(n1673), .CK(clk), .RN(n2239), .Q(
        \register[19][10] ) );
  DFFRX1 \register_reg[19][9]  ( .D(n1674), .CK(clk), .RN(n2239), .Q(
        \register[19][9] ) );
  DFFRX1 \register_reg[23][31]  ( .D(n1780), .CK(clk), .RN(n2231), .Q(
        \register[23][31] ) );
  DFFRX1 \register_reg[23][30]  ( .D(n1781), .CK(clk), .RN(n2231), .Q(
        \register[23][30] ) );
  DFFRX1 \register_reg[23][29]  ( .D(n1782), .CK(clk), .RN(n2230), .Q(
        \register[23][29] ) );
  DFFRX1 \register_reg[23][28]  ( .D(n1783), .CK(clk), .RN(n2230), .Q(
        \register[23][28] ) );
  DFFRX1 \register_reg[23][27]  ( .D(n1784), .CK(clk), .RN(n2230), .Q(
        \register[23][27] ) );
  DFFRX1 \register_reg[23][26]  ( .D(n1785), .CK(clk), .RN(n2230), .Q(
        \register[23][26] ) );
  DFFRX1 \register_reg[23][25]  ( .D(n1786), .CK(clk), .RN(n2230), .Q(
        \register[23][25] ) );
  DFFRX1 \register_reg[23][24]  ( .D(n1787), .CK(clk), .RN(n2230), .Q(
        \register[23][24] ) );
  DFFRX1 \register_reg[23][23]  ( .D(n1788), .CK(clk), .RN(n2230), .Q(
        \register[23][23] ) );
  DFFRX1 \register_reg[23][22]  ( .D(n1789), .CK(clk), .RN(n2230), .Q(
        \register[23][22] ) );
  DFFRX1 \register_reg[23][21]  ( .D(n1790), .CK(clk), .RN(n2230), .Q(
        \register[23][21] ) );
  DFFRX1 \register_reg[23][20]  ( .D(n1791), .CK(clk), .RN(n2230), .Q(
        \register[23][20] ) );
  DFFRX1 \register_reg[23][19]  ( .D(n1792), .CK(clk), .RN(n2230), .Q(
        \register[23][19] ) );
  DFFRX1 \register_reg[23][18]  ( .D(n1793), .CK(clk), .RN(n2230), .Q(
        \register[23][18] ) );
  DFFRX1 \register_reg[23][17]  ( .D(n1794), .CK(clk), .RN(n2230), .Q(
        \register[23][17] ) );
  DFFRX1 \register_reg[23][16]  ( .D(n1795), .CK(clk), .RN(n2229), .Q(
        \register[23][16] ) );
  DFFRX1 \register_reg[23][15]  ( .D(n1796), .CK(clk), .RN(n2229), .Q(
        \register[23][15] ) );
  DFFRX1 \register_reg[23][14]  ( .D(n1797), .CK(clk), .RN(n2229), .Q(
        \register[23][14] ) );
  DFFRX1 \register_reg[23][13]  ( .D(n1798), .CK(clk), .RN(n2229), .Q(
        \register[23][13] ) );
  DFFRX1 \register_reg[23][12]  ( .D(n1799), .CK(clk), .RN(n2229), .Q(
        \register[23][12] ) );
  DFFRX1 \register_reg[23][11]  ( .D(n1800), .CK(clk), .RN(n2229), .Q(
        \register[23][11] ) );
  DFFRX1 \register_reg[23][10]  ( .D(n1801), .CK(clk), .RN(n2229), .Q(
        \register[23][10] ) );
  DFFRX1 \register_reg[23][9]  ( .D(n1802), .CK(clk), .RN(n2229), .Q(
        \register[23][9] ) );
  DFFRX1 \register_reg[27][31]  ( .D(n1908), .CK(clk), .RN(n2221), .Q(
        \register[27][31] ) );
  DFFRX1 \register_reg[27][30]  ( .D(n1909), .CK(clk), .RN(n2221), .Q(
        \register[27][30] ) );
  DFFRX1 \register_reg[27][29]  ( .D(n1910), .CK(clk), .RN(n2221), .Q(
        \register[27][29] ) );
  DFFRX1 \register_reg[27][28]  ( .D(n1911), .CK(clk), .RN(n2221), .Q(
        \register[27][28] ) );
  DFFRX1 \register_reg[27][27]  ( .D(n1912), .CK(clk), .RN(n2220), .Q(
        \register[27][27] ) );
  DFFRX1 \register_reg[27][26]  ( .D(n1913), .CK(clk), .RN(n2220), .Q(
        \register[27][26] ) );
  DFFRX1 \register_reg[27][25]  ( .D(n1914), .CK(clk), .RN(n2220), .Q(
        \register[27][25] ) );
  DFFRX1 \register_reg[27][24]  ( .D(n1915), .CK(clk), .RN(n2220), .Q(
        \register[27][24] ) );
  DFFRX1 \register_reg[27][23]  ( .D(n1916), .CK(clk), .RN(n2220), .Q(
        \register[27][23] ) );
  DFFRX1 \register_reg[27][22]  ( .D(n1917), .CK(clk), .RN(n2220), .Q(
        \register[27][22] ) );
  DFFRX1 \register_reg[27][21]  ( .D(n1918), .CK(clk), .RN(n2220), .Q(
        \register[27][21] ) );
  DFFRX1 \register_reg[27][20]  ( .D(n1919), .CK(clk), .RN(n2220), .Q(
        \register[27][20] ) );
  DFFRX1 \register_reg[27][19]  ( .D(n1920), .CK(clk), .RN(n2220), .Q(
        \register[27][19] ) );
  DFFRX1 \register_reg[27][18]  ( .D(n1921), .CK(clk), .RN(n2220), .Q(
        \register[27][18] ) );
  DFFRX1 \register_reg[27][17]  ( .D(n1922), .CK(clk), .RN(n2220), .Q(
        \register[27][17] ) );
  DFFRX1 \register_reg[27][16]  ( .D(n1923), .CK(clk), .RN(n2220), .Q(
        \register[27][16] ) );
  DFFRX1 \register_reg[27][15]  ( .D(n1924), .CK(clk), .RN(n2220), .Q(
        \register[27][15] ) );
  DFFRX1 \register_reg[27][14]  ( .D(n1925), .CK(clk), .RN(n2219), .Q(
        \register[27][14] ) );
  DFFRX1 \register_reg[27][13]  ( .D(n1926), .CK(clk), .RN(n2219), .Q(
        \register[27][13] ) );
  DFFRX1 \register_reg[27][12]  ( .D(n1927), .CK(clk), .RN(n2219), .Q(
        \register[27][12] ) );
  DFFRX1 \register_reg[27][11]  ( .D(n1928), .CK(clk), .RN(n2219), .Q(
        \register[27][11] ) );
  DFFRX1 \register_reg[27][10]  ( .D(n1929), .CK(clk), .RN(n2219), .Q(
        \register[27][10] ) );
  DFFRX1 \register_reg[27][9]  ( .D(n1930), .CK(clk), .RN(n2219), .Q(
        \register[27][9] ) );
  DFFRX1 \register_reg[31][31]  ( .D(n2036), .CK(clk), .RN(n2211), .Q(
        \register[31][31] ) );
  DFFRX1 \register_reg[31][30]  ( .D(n2037), .CK(clk), .RN(n2211), .Q(
        \register[31][30] ) );
  DFFRX1 \register_reg[31][29]  ( .D(n2038), .CK(clk), .RN(n2211), .Q(
        \register[31][29] ) );
  DFFRX1 \register_reg[31][28]  ( .D(n2039), .CK(clk), .RN(n2211), .Q(
        \register[31][28] ) );
  DFFRX1 \register_reg[31][27]  ( .D(n2040), .CK(clk), .RN(n2211), .Q(
        \register[31][27] ) );
  DFFRX1 \register_reg[31][26]  ( .D(n2041), .CK(clk), .RN(n2211), .Q(
        \register[31][26] ) );
  DFFRX1 \register_reg[31][25]  ( .D(n2042), .CK(clk), .RN(n2210), .Q(
        \register[31][25] ) );
  DFFRX1 \register_reg[31][24]  ( .D(n2043), .CK(clk), .RN(n2210), .Q(
        \register[31][24] ) );
  DFFRX1 \register_reg[31][23]  ( .D(n2044), .CK(clk), .RN(n2210), .Q(
        \register[31][23] ) );
  DFFRX1 \register_reg[31][22]  ( .D(n2045), .CK(clk), .RN(n2210), .Q(
        \register[31][22] ) );
  DFFRX1 \register_reg[31][21]  ( .D(n2046), .CK(clk), .RN(n2210), .Q(
        \register[31][21] ) );
  DFFRX1 \register_reg[31][20]  ( .D(n2047), .CK(clk), .RN(n2210), .Q(
        \register[31][20] ) );
  DFFRX1 \register_reg[31][19]  ( .D(n2048), .CK(clk), .RN(n2210), .Q(
        \register[31][19] ) );
  DFFRX1 \register_reg[31][18]  ( .D(n2049), .CK(clk), .RN(n2210), .Q(
        \register[31][18] ) );
  DFFRX1 \register_reg[31][17]  ( .D(n2050), .CK(clk), .RN(n2210), .Q(
        \register[31][17] ) );
  DFFRX1 \register_reg[31][16]  ( .D(n2051), .CK(clk), .RN(n2210), .Q(
        \register[31][16] ) );
  DFFRX1 \register_reg[31][15]  ( .D(n2052), .CK(clk), .RN(n2210), .Q(
        \register[31][15] ) );
  DFFRX1 \register_reg[31][14]  ( .D(n2053), .CK(clk), .RN(n2210), .Q(
        \register[31][14] ) );
  DFFRX1 \register_reg[31][13]  ( .D(n2054), .CK(clk), .RN(n2210), .Q(
        \register[31][13] ) );
  DFFRX1 \register_reg[31][12]  ( .D(n2055), .CK(clk), .RN(n2209), .Q(
        \register[31][12] ) );
  DFFRX1 \register_reg[31][11]  ( .D(n2056), .CK(clk), .RN(n2209), .Q(
        \register[31][11] ) );
  DFFRX1 \register_reg[31][10]  ( .D(n2057), .CK(clk), .RN(n2209), .Q(
        \register[31][10] ) );
  DFFRX1 \register_reg[31][9]  ( .D(n2058), .CK(clk), .RN(n2209), .Q(
        \register[31][9] ) );
  DFFRX1 \register_reg[1][31]  ( .D(n1076), .CK(clk), .RN(n2285), .Q(
        \register[1][31] ) );
  DFFRX1 \register_reg[1][30]  ( .D(n1077), .CK(clk), .RN(n2285), .Q(
        \register[1][30] ) );
  DFFRX1 \register_reg[1][29]  ( .D(n1078), .CK(clk), .RN(n2285), .Q(
        \register[1][29] ) );
  DFFRX1 \register_reg[1][28]  ( .D(n1079), .CK(clk), .RN(n2285), .Q(
        \register[1][28] ) );
  DFFRX1 \register_reg[1][27]  ( .D(n1080), .CK(clk), .RN(n2284), .Q(
        \register[1][27] ) );
  DFFRX1 \register_reg[1][26]  ( .D(n1081), .CK(clk), .RN(n2284), .Q(
        \register[1][26] ) );
  DFFRX1 \register_reg[1][25]  ( .D(n1082), .CK(clk), .RN(n2284), .Q(
        \register[1][25] ) );
  DFFRX1 \register_reg[1][24]  ( .D(n1083), .CK(clk), .RN(n2284), .Q(
        \register[1][24] ) );
  DFFRX1 \register_reg[1][23]  ( .D(n1084), .CK(clk), .RN(n2284), .Q(
        \register[1][23] ) );
  DFFRX1 \register_reg[1][22]  ( .D(n1085), .CK(clk), .RN(n2284), .Q(
        \register[1][22] ) );
  DFFRX1 \register_reg[1][21]  ( .D(n1086), .CK(clk), .RN(n2284), .Q(
        \register[1][21] ) );
  DFFRX1 \register_reg[1][20]  ( .D(n1087), .CK(clk), .RN(n2284), .Q(
        \register[1][20] ) );
  DFFRX1 \register_reg[1][19]  ( .D(n1088), .CK(clk), .RN(n2284), .Q(
        \register[1][19] ) );
  DFFRX1 \register_reg[1][18]  ( .D(n1089), .CK(clk), .RN(n2284), .Q(
        \register[1][18] ) );
  DFFRX1 \register_reg[1][17]  ( .D(n1090), .CK(clk), .RN(n2284), .Q(
        \register[1][17] ) );
  DFFRX1 \register_reg[1][16]  ( .D(n1091), .CK(clk), .RN(n2284), .Q(
        \register[1][16] ) );
  DFFRX1 \register_reg[1][15]  ( .D(n1092), .CK(clk), .RN(n2284), .Q(
        \register[1][15] ) );
  DFFRX1 \register_reg[1][14]  ( .D(n1093), .CK(clk), .RN(n2283), .Q(
        \register[1][14] ) );
  DFFRX1 \register_reg[1][13]  ( .D(n1094), .CK(clk), .RN(n2283), .Q(
        \register[1][13] ) );
  DFFRX1 \register_reg[1][12]  ( .D(n1095), .CK(clk), .RN(n2283), .Q(
        \register[1][12] ) );
  DFFRX1 \register_reg[1][11]  ( .D(n1096), .CK(clk), .RN(n2283), .Q(
        \register[1][11] ) );
  DFFRX1 \register_reg[1][10]  ( .D(n1097), .CK(clk), .RN(n2283), .Q(
        \register[1][10] ) );
  DFFRX1 \register_reg[1][9]  ( .D(n1098), .CK(clk), .RN(n2283), .Q(
        \register[1][9] ) );
  DFFRX1 \register_reg[5][31]  ( .D(n1204), .CK(clk), .RN(n2275), .Q(
        \register[5][31] ) );
  DFFRX1 \register_reg[5][30]  ( .D(n1205), .CK(clk), .RN(n2275), .Q(
        \register[5][30] ) );
  DFFRX1 \register_reg[5][29]  ( .D(n1206), .CK(clk), .RN(n2275), .Q(
        \register[5][29] ) );
  DFFRX1 \register_reg[5][28]  ( .D(n1207), .CK(clk), .RN(n2275), .Q(
        \register[5][28] ) );
  DFFRX1 \register_reg[5][27]  ( .D(n1208), .CK(clk), .RN(n2275), .Q(
        \register[5][27] ) );
  DFFRX1 \register_reg[5][26]  ( .D(n1209), .CK(clk), .RN(n2275), .Q(
        \register[5][26] ) );
  DFFRX1 \register_reg[5][25]  ( .D(n1210), .CK(clk), .RN(n2274), .Q(
        \register[5][25] ) );
  DFFRX1 \register_reg[5][24]  ( .D(n1211), .CK(clk), .RN(n2274), .Q(
        \register[5][24] ) );
  DFFRX1 \register_reg[5][23]  ( .D(n1212), .CK(clk), .RN(n2274), .Q(
        \register[5][23] ) );
  DFFRX1 \register_reg[5][22]  ( .D(n1213), .CK(clk), .RN(n2274), .Q(
        \register[5][22] ) );
  DFFRX1 \register_reg[5][21]  ( .D(n1214), .CK(clk), .RN(n2274), .Q(
        \register[5][21] ) );
  DFFRX1 \register_reg[5][20]  ( .D(n1215), .CK(clk), .RN(n2274), .Q(
        \register[5][20] ) );
  DFFRX1 \register_reg[5][19]  ( .D(n1216), .CK(clk), .RN(n2274), .Q(
        \register[5][19] ) );
  DFFRX1 \register_reg[5][18]  ( .D(n1217), .CK(clk), .RN(n2274), .Q(
        \register[5][18] ) );
  DFFRX1 \register_reg[5][17]  ( .D(n1218), .CK(clk), .RN(n2274), .Q(
        \register[5][17] ) );
  DFFRX1 \register_reg[5][16]  ( .D(n1219), .CK(clk), .RN(n2274), .Q(
        \register[5][16] ) );
  DFFRX1 \register_reg[5][15]  ( .D(n1220), .CK(clk), .RN(n2274), .Q(
        \register[5][15] ) );
  DFFRX1 \register_reg[5][14]  ( .D(n1221), .CK(clk), .RN(n2274), .Q(
        \register[5][14] ) );
  DFFRX1 \register_reg[5][13]  ( .D(n1222), .CK(clk), .RN(n2274), .Q(
        \register[5][13] ) );
  DFFRX1 \register_reg[5][12]  ( .D(n1223), .CK(clk), .RN(n2273), .Q(
        \register[5][12] ) );
  DFFRX1 \register_reg[5][11]  ( .D(n1224), .CK(clk), .RN(n2273), .Q(
        \register[5][11] ) );
  DFFRX1 \register_reg[5][10]  ( .D(n1225), .CK(clk), .RN(n2273), .Q(
        \register[5][10] ) );
  DFFRX1 \register_reg[5][9]  ( .D(n1226), .CK(clk), .RN(n2273), .Q(
        \register[5][9] ) );
  DFFRX1 \register_reg[9][31]  ( .D(n1332), .CK(clk), .RN(n2265), .Q(
        \register[9][31] ) );
  DFFRX1 \register_reg[9][30]  ( .D(n1333), .CK(clk), .RN(n2265), .Q(
        \register[9][30] ) );
  DFFRX1 \register_reg[9][29]  ( .D(n1334), .CK(clk), .RN(n2265), .Q(
        \register[9][29] ) );
  DFFRX1 \register_reg[9][28]  ( .D(n1335), .CK(clk), .RN(n2265), .Q(
        \register[9][28] ) );
  DFFRX1 \register_reg[9][27]  ( .D(n1336), .CK(clk), .RN(n2265), .Q(
        \register[9][27] ) );
  DFFRX1 \register_reg[9][26]  ( .D(n1337), .CK(clk), .RN(n2265), .Q(
        \register[9][26] ) );
  DFFRX1 \register_reg[9][25]  ( .D(n1338), .CK(clk), .RN(n2265), .Q(
        \register[9][25] ) );
  DFFRX1 \register_reg[9][24]  ( .D(n1339), .CK(clk), .RN(n2265), .Q(
        \register[9][24] ) );
  DFFRX1 \register_reg[9][23]  ( .D(n1340), .CK(clk), .RN(n2264), .Q(
        \register[9][23] ) );
  DFFRX1 \register_reg[9][22]  ( .D(n1341), .CK(clk), .RN(n2264), .Q(
        \register[9][22] ) );
  DFFRX1 \register_reg[9][21]  ( .D(n1342), .CK(clk), .RN(n2264), .Q(
        \register[9][21] ) );
  DFFRX1 \register_reg[9][20]  ( .D(n1343), .CK(clk), .RN(n2264), .Q(
        \register[9][20] ) );
  DFFRX1 \register_reg[9][19]  ( .D(n1344), .CK(clk), .RN(n2264), .Q(
        \register[9][19] ) );
  DFFRX1 \register_reg[9][18]  ( .D(n1345), .CK(clk), .RN(n2264), .Q(
        \register[9][18] ) );
  DFFRX1 \register_reg[9][17]  ( .D(n1346), .CK(clk), .RN(n2264), .Q(
        \register[9][17] ) );
  DFFRX1 \register_reg[9][16]  ( .D(n1347), .CK(clk), .RN(n2264), .Q(
        \register[9][16] ) );
  DFFRX1 \register_reg[9][15]  ( .D(n1348), .CK(clk), .RN(n2264), .Q(
        \register[9][15] ) );
  DFFRX1 \register_reg[9][14]  ( .D(n1349), .CK(clk), .RN(n2264), .Q(
        \register[9][14] ) );
  DFFRX1 \register_reg[9][13]  ( .D(n1350), .CK(clk), .RN(n2264), .Q(
        \register[9][13] ) );
  DFFRX1 \register_reg[9][12]  ( .D(n1351), .CK(clk), .RN(n2264), .Q(
        \register[9][12] ) );
  DFFRX1 \register_reg[9][11]  ( .D(n1352), .CK(clk), .RN(n2264), .Q(
        \register[9][11] ) );
  DFFRX1 \register_reg[9][10]  ( .D(n1353), .CK(clk), .RN(n2263), .Q(
        \register[9][10] ) );
  DFFRX1 \register_reg[9][9]  ( .D(n1354), .CK(clk), .RN(n2263), .Q(
        \register[9][9] ) );
  DFFRX1 \register_reg[13][31]  ( .D(n1460), .CK(clk), .RN(n2255), .Q(
        \register[13][31] ) );
  DFFRX1 \register_reg[13][30]  ( .D(n1461), .CK(clk), .RN(n2255), .Q(
        \register[13][30] ) );
  DFFRX1 \register_reg[13][29]  ( .D(n1462), .CK(clk), .RN(n2255), .Q(
        \register[13][29] ) );
  DFFRX1 \register_reg[13][28]  ( .D(n1463), .CK(clk), .RN(n2255), .Q(
        \register[13][28] ) );
  DFFRX1 \register_reg[13][27]  ( .D(n1464), .CK(clk), .RN(n2255), .Q(
        \register[13][27] ) );
  DFFRX1 \register_reg[13][26]  ( .D(n1465), .CK(clk), .RN(n2255), .Q(
        \register[13][26] ) );
  DFFRX1 \register_reg[13][25]  ( .D(n1466), .CK(clk), .RN(n2255), .Q(
        \register[13][25] ) );
  DFFRX1 \register_reg[13][24]  ( .D(n1467), .CK(clk), .RN(n2255), .Q(
        \register[13][24] ) );
  DFFRX1 \register_reg[13][23]  ( .D(n1468), .CK(clk), .RN(n2255), .Q(
        \register[13][23] ) );
  DFFRX1 \register_reg[13][22]  ( .D(n1469), .CK(clk), .RN(n2255), .Q(
        \register[13][22] ) );
  DFFRX1 \register_reg[13][21]  ( .D(n1470), .CK(clk), .RN(n2254), .Q(
        \register[13][21] ) );
  DFFRX1 \register_reg[13][20]  ( .D(n1471), .CK(clk), .RN(n2254), .Q(
        \register[13][20] ) );
  DFFRX1 \register_reg[13][19]  ( .D(n1472), .CK(clk), .RN(n2254), .Q(
        \register[13][19] ) );
  DFFRX1 \register_reg[13][18]  ( .D(n1473), .CK(clk), .RN(n2254), .Q(
        \register[13][18] ) );
  DFFRX1 \register_reg[13][17]  ( .D(n1474), .CK(clk), .RN(n2254), .Q(
        \register[13][17] ) );
  DFFRX1 \register_reg[13][16]  ( .D(n1475), .CK(clk), .RN(n2254), .Q(
        \register[13][16] ) );
  DFFRX1 \register_reg[13][15]  ( .D(n1476), .CK(clk), .RN(n2254), .Q(
        \register[13][15] ) );
  DFFRX1 \register_reg[13][14]  ( .D(n1477), .CK(clk), .RN(n2254), .Q(
        \register[13][14] ) );
  DFFRX1 \register_reg[13][13]  ( .D(n1478), .CK(clk), .RN(n2254), .Q(
        \register[13][13] ) );
  DFFRX1 \register_reg[13][12]  ( .D(n1479), .CK(clk), .RN(n2254), .Q(
        \register[13][12] ) );
  DFFRX1 \register_reg[13][11]  ( .D(n1480), .CK(clk), .RN(n2254), .Q(
        \register[13][11] ) );
  DFFRX1 \register_reg[13][10]  ( .D(n1481), .CK(clk), .RN(n2254), .Q(
        \register[13][10] ) );
  DFFRX1 \register_reg[13][9]  ( .D(n1482), .CK(clk), .RN(n2254), .Q(
        \register[13][9] ) );
  DFFRX1 \register_reg[17][31]  ( .D(n1588), .CK(clk), .RN(n2245), .Q(
        \register[17][31] ) );
  DFFRX1 \register_reg[17][30]  ( .D(n1589), .CK(clk), .RN(n2245), .Q(
        \register[17][30] ) );
  DFFRX1 \register_reg[17][29]  ( .D(n1590), .CK(clk), .RN(n2245), .Q(
        \register[17][29] ) );
  DFFRX1 \register_reg[17][28]  ( .D(n1591), .CK(clk), .RN(n2245), .Q(
        \register[17][28] ) );
  DFFRX1 \register_reg[17][27]  ( .D(n1592), .CK(clk), .RN(n2245), .Q(
        \register[17][27] ) );
  DFFRX1 \register_reg[17][26]  ( .D(n1593), .CK(clk), .RN(n2245), .Q(
        \register[17][26] ) );
  DFFRX1 \register_reg[17][25]  ( .D(n1594), .CK(clk), .RN(n2245), .Q(
        \register[17][25] ) );
  DFFRX1 \register_reg[17][24]  ( .D(n1595), .CK(clk), .RN(n2245), .Q(
        \register[17][24] ) );
  DFFRX1 \register_reg[17][23]  ( .D(n1596), .CK(clk), .RN(n2245), .Q(
        \register[17][23] ) );
  DFFRX1 \register_reg[17][22]  ( .D(n1597), .CK(clk), .RN(n2245), .Q(
        \register[17][22] ) );
  DFFRX1 \register_reg[17][21]  ( .D(n1598), .CK(clk), .RN(n2245), .Q(
        \register[17][21] ) );
  DFFRX1 \register_reg[17][20]  ( .D(n1599), .CK(clk), .RN(n2245), .Q(
        \register[17][20] ) );
  DFFRX1 \register_reg[17][19]  ( .D(n1600), .CK(clk), .RN(n2244), .Q(
        \register[17][19] ) );
  DFFRX1 \register_reg[17][18]  ( .D(n1601), .CK(clk), .RN(n2244), .Q(
        \register[17][18] ) );
  DFFRX1 \register_reg[17][17]  ( .D(n1602), .CK(clk), .RN(n2244), .Q(
        \register[17][17] ) );
  DFFRX1 \register_reg[17][16]  ( .D(n1603), .CK(clk), .RN(n2244), .Q(
        \register[17][16] ) );
  DFFRX1 \register_reg[17][15]  ( .D(n1604), .CK(clk), .RN(n2244), .Q(
        \register[17][15] ) );
  DFFRX1 \register_reg[17][14]  ( .D(n1605), .CK(clk), .RN(n2244), .Q(
        \register[17][14] ) );
  DFFRX1 \register_reg[17][13]  ( .D(n1606), .CK(clk), .RN(n2244), .Q(
        \register[17][13] ) );
  DFFRX1 \register_reg[17][12]  ( .D(n1607), .CK(clk), .RN(n2244), .Q(
        \register[17][12] ) );
  DFFRX1 \register_reg[17][11]  ( .D(n1608), .CK(clk), .RN(n2244), .Q(
        \register[17][11] ) );
  DFFRX1 \register_reg[17][10]  ( .D(n1609), .CK(clk), .RN(n2244), .Q(
        \register[17][10] ) );
  DFFRX1 \register_reg[17][9]  ( .D(n1610), .CK(clk), .RN(n2244), .Q(
        \register[17][9] ) );
  DFFRX1 \register_reg[21][31]  ( .D(n1716), .CK(clk), .RN(n2236), .Q(
        \register[21][31] ) );
  DFFRX1 \register_reg[21][30]  ( .D(n1717), .CK(clk), .RN(n2235), .Q(
        \register[21][30] ) );
  DFFRX1 \register_reg[21][29]  ( .D(n1718), .CK(clk), .RN(n2235), .Q(
        \register[21][29] ) );
  DFFRX1 \register_reg[21][28]  ( .D(n1719), .CK(clk), .RN(n2235), .Q(
        \register[21][28] ) );
  DFFRX1 \register_reg[21][27]  ( .D(n1720), .CK(clk), .RN(n2235), .Q(
        \register[21][27] ) );
  DFFRX1 \register_reg[21][26]  ( .D(n1721), .CK(clk), .RN(n2235), .Q(
        \register[21][26] ) );
  DFFRX1 \register_reg[21][25]  ( .D(n1722), .CK(clk), .RN(n2235), .Q(
        \register[21][25] ) );
  DFFRX1 \register_reg[21][24]  ( .D(n1723), .CK(clk), .RN(n2235), .Q(
        \register[21][24] ) );
  DFFRX1 \register_reg[21][23]  ( .D(n1724), .CK(clk), .RN(n2235), .Q(
        \register[21][23] ) );
  DFFRX1 \register_reg[21][22]  ( .D(n1725), .CK(clk), .RN(n2235), .Q(
        \register[21][22] ) );
  DFFRX1 \register_reg[21][21]  ( .D(n1726), .CK(clk), .RN(n2235), .Q(
        \register[21][21] ) );
  DFFRX1 \register_reg[21][20]  ( .D(n1727), .CK(clk), .RN(n2235), .Q(
        \register[21][20] ) );
  DFFRX1 \register_reg[21][19]  ( .D(n1728), .CK(clk), .RN(n2235), .Q(
        \register[21][19] ) );
  DFFRX1 \register_reg[21][18]  ( .D(n1729), .CK(clk), .RN(n2235), .Q(
        \register[21][18] ) );
  DFFRX1 \register_reg[21][17]  ( .D(n1730), .CK(clk), .RN(n2234), .Q(
        \register[21][17] ) );
  DFFRX1 \register_reg[21][16]  ( .D(n1731), .CK(clk), .RN(n2234), .Q(
        \register[21][16] ) );
  DFFRX1 \register_reg[21][15]  ( .D(n1732), .CK(clk), .RN(n2234), .Q(
        \register[21][15] ) );
  DFFRX1 \register_reg[21][14]  ( .D(n1733), .CK(clk), .RN(n2234), .Q(
        \register[21][14] ) );
  DFFRX1 \register_reg[21][13]  ( .D(n1734), .CK(clk), .RN(n2234), .Q(
        \register[21][13] ) );
  DFFRX1 \register_reg[21][12]  ( .D(n1735), .CK(clk), .RN(n2234), .Q(
        \register[21][12] ) );
  DFFRX1 \register_reg[21][11]  ( .D(n1736), .CK(clk), .RN(n2234), .Q(
        \register[21][11] ) );
  DFFRX1 \register_reg[21][10]  ( .D(n1737), .CK(clk), .RN(n2234), .Q(
        \register[21][10] ) );
  DFFRX1 \register_reg[21][9]  ( .D(n1738), .CK(clk), .RN(n2234), .Q(
        \register[21][9] ) );
  DFFRX1 \register_reg[25][31]  ( .D(n1844), .CK(clk), .RN(n2226), .Q(
        \register[25][31] ) );
  DFFRX1 \register_reg[25][30]  ( .D(n1845), .CK(clk), .RN(n2226), .Q(
        \register[25][30] ) );
  DFFRX1 \register_reg[25][29]  ( .D(n1846), .CK(clk), .RN(n2226), .Q(
        \register[25][29] ) );
  DFFRX1 \register_reg[25][28]  ( .D(n1847), .CK(clk), .RN(n2225), .Q(
        \register[25][28] ) );
  DFFRX1 \register_reg[25][27]  ( .D(n1848), .CK(clk), .RN(n2225), .Q(
        \register[25][27] ) );
  DFFRX1 \register_reg[25][26]  ( .D(n1849), .CK(clk), .RN(n2225), .Q(
        \register[25][26] ) );
  DFFRX1 \register_reg[25][25]  ( .D(n1850), .CK(clk), .RN(n2225), .Q(
        \register[25][25] ) );
  DFFRX1 \register_reg[25][24]  ( .D(n1851), .CK(clk), .RN(n2225), .Q(
        \register[25][24] ) );
  DFFRX1 \register_reg[25][23]  ( .D(n1852), .CK(clk), .RN(n2225), .Q(
        \register[25][23] ) );
  DFFRX1 \register_reg[25][22]  ( .D(n1853), .CK(clk), .RN(n2225), .Q(
        \register[25][22] ) );
  DFFRX1 \register_reg[25][21]  ( .D(n1854), .CK(clk), .RN(n2225), .Q(
        \register[25][21] ) );
  DFFRX1 \register_reg[25][20]  ( .D(n1855), .CK(clk), .RN(n2225), .Q(
        \register[25][20] ) );
  DFFRX1 \register_reg[25][19]  ( .D(n1856), .CK(clk), .RN(n2225), .Q(
        \register[25][19] ) );
  DFFRX1 \register_reg[25][18]  ( .D(n1857), .CK(clk), .RN(n2225), .Q(
        \register[25][18] ) );
  DFFRX1 \register_reg[25][17]  ( .D(n1858), .CK(clk), .RN(n2225), .Q(
        \register[25][17] ) );
  DFFRX1 \register_reg[25][16]  ( .D(n1859), .CK(clk), .RN(n2225), .Q(
        \register[25][16] ) );
  DFFRX1 \register_reg[25][15]  ( .D(n1860), .CK(clk), .RN(n2224), .Q(
        \register[25][15] ) );
  DFFRX1 \register_reg[25][14]  ( .D(n1861), .CK(clk), .RN(n2224), .Q(
        \register[25][14] ) );
  DFFRX1 \register_reg[25][13]  ( .D(n1862), .CK(clk), .RN(n2224), .Q(
        \register[25][13] ) );
  DFFRX1 \register_reg[25][12]  ( .D(n1863), .CK(clk), .RN(n2224), .Q(
        \register[25][12] ) );
  DFFRX1 \register_reg[25][11]  ( .D(n1864), .CK(clk), .RN(n2224), .Q(
        \register[25][11] ) );
  DFFRX1 \register_reg[25][10]  ( .D(n1865), .CK(clk), .RN(n2224), .Q(
        \register[25][10] ) );
  DFFRX1 \register_reg[25][9]  ( .D(n1866), .CK(clk), .RN(n2224), .Q(
        \register[25][9] ) );
  DFFRX1 \register_reg[29][31]  ( .D(n1972), .CK(clk), .RN(n2216), .Q(
        \register[29][31] ) );
  DFFRX1 \register_reg[29][30]  ( .D(n1973), .CK(clk), .RN(n2216), .Q(
        \register[29][30] ) );
  DFFRX1 \register_reg[29][29]  ( .D(n1974), .CK(clk), .RN(n2216), .Q(
        \register[29][29] ) );
  DFFRX1 \register_reg[29][28]  ( .D(n1975), .CK(clk), .RN(n2216), .Q(
        \register[29][28] ) );
  DFFRX1 \register_reg[29][27]  ( .D(n1976), .CK(clk), .RN(n2216), .Q(
        \register[29][27] ) );
  DFFRX1 \register_reg[29][26]  ( .D(n1977), .CK(clk), .RN(n2215), .Q(
        \register[29][26] ) );
  DFFRX1 \register_reg[29][25]  ( .D(n1978), .CK(clk), .RN(n2215), .Q(
        \register[29][25] ) );
  DFFRX1 \register_reg[29][24]  ( .D(n1979), .CK(clk), .RN(n2215), .Q(
        \register[29][24] ) );
  DFFRX1 \register_reg[29][23]  ( .D(n1980), .CK(clk), .RN(n2215), .Q(
        \register[29][23] ) );
  DFFRX1 \register_reg[29][22]  ( .D(n1981), .CK(clk), .RN(n2215), .Q(
        \register[29][22] ) );
  DFFRX1 \register_reg[29][21]  ( .D(n1982), .CK(clk), .RN(n2215), .Q(
        \register[29][21] ) );
  DFFRX1 \register_reg[29][20]  ( .D(n1983), .CK(clk), .RN(n2215), .Q(
        \register[29][20] ) );
  DFFRX1 \register_reg[29][19]  ( .D(n1984), .CK(clk), .RN(n2215), .Q(
        \register[29][19] ) );
  DFFRX1 \register_reg[29][18]  ( .D(n1985), .CK(clk), .RN(n2215), .Q(
        \register[29][18] ) );
  DFFRX1 \register_reg[29][17]  ( .D(n1986), .CK(clk), .RN(n2215), .Q(
        \register[29][17] ) );
  DFFRX1 \register_reg[29][16]  ( .D(n1987), .CK(clk), .RN(n2215), .Q(
        \register[29][16] ) );
  DFFRX1 \register_reg[29][15]  ( .D(n1988), .CK(clk), .RN(n2215), .Q(
        \register[29][15] ) );
  DFFRX1 \register_reg[29][14]  ( .D(n1989), .CK(clk), .RN(n2215), .Q(
        \register[29][14] ) );
  DFFRX1 \register_reg[29][13]  ( .D(n1990), .CK(clk), .RN(n2214), .Q(
        \register[29][13] ) );
  DFFRX1 \register_reg[29][12]  ( .D(n1991), .CK(clk), .RN(n2214), .Q(
        \register[29][12] ) );
  DFFRX1 \register_reg[29][11]  ( .D(n1992), .CK(clk), .RN(n2214), .Q(
        \register[29][11] ) );
  DFFRX1 \register_reg[29][10]  ( .D(n1993), .CK(clk), .RN(n2214), .Q(
        \register[29][10] ) );
  DFFRX1 \register_reg[29][9]  ( .D(n1994), .CK(clk), .RN(n2214), .Q(
        \register[29][9] ) );
  DFFRX1 \register_reg[0][31]  ( .D(n1044), .CK(clk), .RN(n2287), .Q(
        \register[0][31] ) );
  DFFRX1 \register_reg[0][30]  ( .D(n1045), .CK(clk), .RN(n2287), .Q(
        \register[0][30] ) );
  DFFRX1 \register_reg[0][29]  ( .D(n1046), .CK(clk), .RN(n2287), .Q(
        \register[0][29] ) );
  DFFRX1 \register_reg[0][28]  ( .D(n1047), .CK(clk), .RN(n2287), .Q(
        \register[0][28] ) );
  DFFRX1 \register_reg[0][27]  ( .D(n1048), .CK(clk), .RN(n2287), .Q(
        \register[0][27] ) );
  DFFRX1 \register_reg[0][26]  ( .D(n1049), .CK(clk), .RN(n2287), .Q(
        \register[0][26] ) );
  DFFRX1 \register_reg[0][25]  ( .D(n1050), .CK(clk), .RN(n2287), .Q(
        \register[0][25] ) );
  DFFRX1 \register_reg[0][24]  ( .D(n1051), .CK(clk), .RN(n2287), .Q(
        \register[0][24] ) );
  DFFRX1 \register_reg[0][23]  ( .D(n1052), .CK(clk), .RN(n2287), .Q(
        \register[0][23] ) );
  DFFRX1 \register_reg[0][22]  ( .D(n1053), .CK(clk), .RN(n2287), .Q(
        \register[0][22] ) );
  DFFRX1 \register_reg[0][21]  ( .D(n1054), .CK(clk), .RN(n2286), .Q(
        \register[0][21] ) );
  DFFRX1 \register_reg[0][20]  ( .D(n1055), .CK(clk), .RN(n2286), .Q(
        \register[0][20] ) );
  DFFRX1 \register_reg[0][19]  ( .D(n1056), .CK(clk), .RN(n2286), .Q(
        \register[0][19] ) );
  DFFRX1 \register_reg[0][18]  ( .D(n1057), .CK(clk), .RN(n2286), .Q(
        \register[0][18] ) );
  DFFRX1 \register_reg[0][17]  ( .D(n1058), .CK(clk), .RN(n2286), .Q(
        \register[0][17] ) );
  DFFRX1 \register_reg[0][16]  ( .D(n1059), .CK(clk), .RN(n2286), .Q(
        \register[0][16] ) );
  DFFRX1 \register_reg[0][15]  ( .D(n1060), .CK(clk), .RN(n2286), .Q(
        \register[0][15] ) );
  DFFRX1 \register_reg[0][14]  ( .D(n1061), .CK(clk), .RN(n2286), .Q(
        \register[0][14] ) );
  DFFRX1 \register_reg[0][13]  ( .D(n1062), .CK(clk), .RN(n2286), .Q(
        \register[0][13] ) );
  DFFRX1 \register_reg[0][12]  ( .D(n1063), .CK(clk), .RN(n2286), .Q(
        \register[0][12] ) );
  DFFRX1 \register_reg[0][11]  ( .D(n1064), .CK(clk), .RN(n2286), .Q(
        \register[0][11] ) );
  DFFRX1 \register_reg[0][10]  ( .D(n1065), .CK(clk), .RN(n2286), .Q(
        \register[0][10] ) );
  DFFRX1 \register_reg[0][9]  ( .D(n1066), .CK(clk), .RN(n2286), .Q(
        \register[0][9] ) );
  DFFRX1 \register_reg[4][31]  ( .D(n1172), .CK(clk), .RN(n2277), .Q(
        \register[4][31] ) );
  DFFRX1 \register_reg[4][30]  ( .D(n1173), .CK(clk), .RN(n2277), .Q(
        \register[4][30] ) );
  DFFRX1 \register_reg[4][29]  ( .D(n1174), .CK(clk), .RN(n2277), .Q(
        \register[4][29] ) );
  DFFRX1 \register_reg[4][28]  ( .D(n1175), .CK(clk), .RN(n2277), .Q(
        \register[4][28] ) );
  DFFRX1 \register_reg[4][27]  ( .D(n1176), .CK(clk), .RN(n2277), .Q(
        \register[4][27] ) );
  DFFRX1 \register_reg[4][26]  ( .D(n1177), .CK(clk), .RN(n2277), .Q(
        \register[4][26] ) );
  DFFRX1 \register_reg[4][25]  ( .D(n1178), .CK(clk), .RN(n2277), .Q(
        \register[4][25] ) );
  DFFRX1 \register_reg[4][24]  ( .D(n1179), .CK(clk), .RN(n2277), .Q(
        \register[4][24] ) );
  DFFRX1 \register_reg[4][23]  ( .D(n1180), .CK(clk), .RN(n2277), .Q(
        \register[4][23] ) );
  DFFRX1 \register_reg[4][22]  ( .D(n1181), .CK(clk), .RN(n2277), .Q(
        \register[4][22] ) );
  DFFRX1 \register_reg[4][21]  ( .D(n1182), .CK(clk), .RN(n2277), .Q(
        \register[4][21] ) );
  DFFRX1 \register_reg[4][20]  ( .D(n1183), .CK(clk), .RN(n2277), .Q(
        \register[4][20] ) );
  DFFRX1 \register_reg[4][19]  ( .D(n1184), .CK(clk), .RN(n2276), .Q(
        \register[4][19] ) );
  DFFRX1 \register_reg[4][18]  ( .D(n1185), .CK(clk), .RN(n2276), .Q(
        \register[4][18] ) );
  DFFRX1 \register_reg[4][17]  ( .D(n1186), .CK(clk), .RN(n2276), .Q(
        \register[4][17] ) );
  DFFRX1 \register_reg[4][16]  ( .D(n1187), .CK(clk), .RN(n2276), .Q(
        \register[4][16] ) );
  DFFRX1 \register_reg[4][15]  ( .D(n1188), .CK(clk), .RN(n2276), .Q(
        \register[4][15] ) );
  DFFRX1 \register_reg[4][14]  ( .D(n1189), .CK(clk), .RN(n2276), .Q(
        \register[4][14] ) );
  DFFRX1 \register_reg[4][13]  ( .D(n1190), .CK(clk), .RN(n2276), .Q(
        \register[4][13] ) );
  DFFRX1 \register_reg[4][12]  ( .D(n1191), .CK(clk), .RN(n2276), .Q(
        \register[4][12] ) );
  DFFRX1 \register_reg[4][11]  ( .D(n1192), .CK(clk), .RN(n2276), .Q(
        \register[4][11] ) );
  DFFRX1 \register_reg[4][10]  ( .D(n1193), .CK(clk), .RN(n2276), .Q(
        \register[4][10] ) );
  DFFRX1 \register_reg[4][9]  ( .D(n1194), .CK(clk), .RN(n2276), .Q(
        \register[4][9] ) );
  DFFRX1 \register_reg[8][31]  ( .D(n1300), .CK(clk), .RN(n2268), .Q(
        \register[8][31] ) );
  DFFRX1 \register_reg[8][30]  ( .D(n1301), .CK(clk), .RN(n2267), .Q(
        \register[8][30] ) );
  DFFRX1 \register_reg[8][29]  ( .D(n1302), .CK(clk), .RN(n2267), .Q(
        \register[8][29] ) );
  DFFRX1 \register_reg[8][28]  ( .D(n1303), .CK(clk), .RN(n2267), .Q(
        \register[8][28] ) );
  DFFRX1 \register_reg[8][27]  ( .D(n1304), .CK(clk), .RN(n2267), .Q(
        \register[8][27] ) );
  DFFRX1 \register_reg[8][26]  ( .D(n1305), .CK(clk), .RN(n2267), .Q(
        \register[8][26] ) );
  DFFRX1 \register_reg[8][25]  ( .D(n1306), .CK(clk), .RN(n2267), .Q(
        \register[8][25] ) );
  DFFRX1 \register_reg[8][24]  ( .D(n1307), .CK(clk), .RN(n2267), .Q(
        \register[8][24] ) );
  DFFRX1 \register_reg[8][23]  ( .D(n1308), .CK(clk), .RN(n2267), .Q(
        \register[8][23] ) );
  DFFRX1 \register_reg[8][22]  ( .D(n1309), .CK(clk), .RN(n2267), .Q(
        \register[8][22] ) );
  DFFRX1 \register_reg[8][21]  ( .D(n1310), .CK(clk), .RN(n2267), .Q(
        \register[8][21] ) );
  DFFRX1 \register_reg[8][20]  ( .D(n1311), .CK(clk), .RN(n2267), .Q(
        \register[8][20] ) );
  DFFRX1 \register_reg[8][19]  ( .D(n1312), .CK(clk), .RN(n2267), .Q(
        \register[8][19] ) );
  DFFRX1 \register_reg[8][18]  ( .D(n1313), .CK(clk), .RN(n2267), .Q(
        \register[8][18] ) );
  DFFRX1 \register_reg[8][17]  ( .D(n1314), .CK(clk), .RN(n2266), .Q(
        \register[8][17] ) );
  DFFRX1 \register_reg[8][16]  ( .D(n1315), .CK(clk), .RN(n2266), .Q(
        \register[8][16] ) );
  DFFRX1 \register_reg[8][15]  ( .D(n1316), .CK(clk), .RN(n2266), .Q(
        \register[8][15] ) );
  DFFRX1 \register_reg[8][14]  ( .D(n1317), .CK(clk), .RN(n2266), .Q(
        \register[8][14] ) );
  DFFRX1 \register_reg[8][13]  ( .D(n1318), .CK(clk), .RN(n2266), .Q(
        \register[8][13] ) );
  DFFRX1 \register_reg[8][12]  ( .D(n1319), .CK(clk), .RN(n2266), .Q(
        \register[8][12] ) );
  DFFRX1 \register_reg[8][11]  ( .D(n1320), .CK(clk), .RN(n2266), .Q(
        \register[8][11] ) );
  DFFRX1 \register_reg[8][10]  ( .D(n1321), .CK(clk), .RN(n2266), .Q(
        \register[8][10] ) );
  DFFRX1 \register_reg[8][9]  ( .D(n1322), .CK(clk), .RN(n2266), .Q(
        \register[8][9] ) );
  DFFRX1 \register_reg[12][31]  ( .D(n1428), .CK(clk), .RN(n2258), .Q(
        \register[12][31] ) );
  DFFRX1 \register_reg[12][30]  ( .D(n1429), .CK(clk), .RN(n2258), .Q(
        \register[12][30] ) );
  DFFRX1 \register_reg[12][29]  ( .D(n1430), .CK(clk), .RN(n2258), .Q(
        \register[12][29] ) );
  DFFRX1 \register_reg[12][28]  ( .D(n1431), .CK(clk), .RN(n2257), .Q(
        \register[12][28] ) );
  DFFRX1 \register_reg[12][27]  ( .D(n1432), .CK(clk), .RN(n2257), .Q(
        \register[12][27] ) );
  DFFRX1 \register_reg[12][26]  ( .D(n1433), .CK(clk), .RN(n2257), .Q(
        \register[12][26] ) );
  DFFRX1 \register_reg[12][25]  ( .D(n1434), .CK(clk), .RN(n2257), .Q(
        \register[12][25] ) );
  DFFRX1 \register_reg[12][24]  ( .D(n1435), .CK(clk), .RN(n2257), .Q(
        \register[12][24] ) );
  DFFRX1 \register_reg[12][23]  ( .D(n1436), .CK(clk), .RN(n2257), .Q(
        \register[12][23] ) );
  DFFRX1 \register_reg[12][22]  ( .D(n1437), .CK(clk), .RN(n2257), .Q(
        \register[12][22] ) );
  DFFRX1 \register_reg[12][21]  ( .D(n1438), .CK(clk), .RN(n2257), .Q(
        \register[12][21] ) );
  DFFRX1 \register_reg[12][20]  ( .D(n1439), .CK(clk), .RN(n2257), .Q(
        \register[12][20] ) );
  DFFRX1 \register_reg[12][19]  ( .D(n1440), .CK(clk), .RN(n2257), .Q(
        \register[12][19] ) );
  DFFRX1 \register_reg[12][18]  ( .D(n1441), .CK(clk), .RN(n2257), .Q(
        \register[12][18] ) );
  DFFRX1 \register_reg[12][17]  ( .D(n1442), .CK(clk), .RN(n2257), .Q(
        \register[12][17] ) );
  DFFRX1 \register_reg[12][16]  ( .D(n1443), .CK(clk), .RN(n2257), .Q(
        \register[12][16] ) );
  DFFRX1 \register_reg[12][15]  ( .D(n1444), .CK(clk), .RN(n2256), .Q(
        \register[12][15] ) );
  DFFRX1 \register_reg[12][14]  ( .D(n1445), .CK(clk), .RN(n2256), .Q(
        \register[12][14] ) );
  DFFRX1 \register_reg[12][13]  ( .D(n1446), .CK(clk), .RN(n2256), .Q(
        \register[12][13] ) );
  DFFRX1 \register_reg[12][12]  ( .D(n1447), .CK(clk), .RN(n2256), .Q(
        \register[12][12] ) );
  DFFRX1 \register_reg[12][11]  ( .D(n1448), .CK(clk), .RN(n2256), .Q(
        \register[12][11] ) );
  DFFRX1 \register_reg[12][10]  ( .D(n1449), .CK(clk), .RN(n2256), .Q(
        \register[12][10] ) );
  DFFRX1 \register_reg[12][9]  ( .D(n1450), .CK(clk), .RN(n2256), .Q(
        \register[12][9] ) );
  DFFRX1 \register_reg[16][31]  ( .D(n1556), .CK(clk), .RN(n2248), .Q(
        \register[16][31] ) );
  DFFRX1 \register_reg[16][30]  ( .D(n1557), .CK(clk), .RN(n2248), .Q(
        \register[16][30] ) );
  DFFRX1 \register_reg[16][29]  ( .D(n1558), .CK(clk), .RN(n2248), .Q(
        \register[16][29] ) );
  DFFRX1 \register_reg[16][28]  ( .D(n1559), .CK(clk), .RN(n2248), .Q(
        \register[16][28] ) );
  DFFRX1 \register_reg[16][27]  ( .D(n1560), .CK(clk), .RN(n2248), .Q(
        \register[16][27] ) );
  DFFRX1 \register_reg[16][26]  ( .D(n1561), .CK(clk), .RN(n2247), .Q(
        \register[16][26] ) );
  DFFRX1 \register_reg[16][25]  ( .D(n1562), .CK(clk), .RN(n2247), .Q(
        \register[16][25] ) );
  DFFRX1 \register_reg[16][24]  ( .D(n1563), .CK(clk), .RN(n2247), .Q(
        \register[16][24] ) );
  DFFRX1 \register_reg[16][23]  ( .D(n1564), .CK(clk), .RN(n2247), .Q(
        \register[16][23] ) );
  DFFRX1 \register_reg[16][22]  ( .D(n1565), .CK(clk), .RN(n2247), .Q(
        \register[16][22] ) );
  DFFRX1 \register_reg[16][21]  ( .D(n1566), .CK(clk), .RN(n2247), .Q(
        \register[16][21] ) );
  DFFRX1 \register_reg[16][20]  ( .D(n1567), .CK(clk), .RN(n2247), .Q(
        \register[16][20] ) );
  DFFRX1 \register_reg[16][19]  ( .D(n1568), .CK(clk), .RN(n2247), .Q(
        \register[16][19] ) );
  DFFRX1 \register_reg[16][18]  ( .D(n1569), .CK(clk), .RN(n2247), .Q(
        \register[16][18] ) );
  DFFRX1 \register_reg[16][17]  ( .D(n1570), .CK(clk), .RN(n2247), .Q(
        \register[16][17] ) );
  DFFRX1 \register_reg[16][16]  ( .D(n1571), .CK(clk), .RN(n2247), .Q(
        \register[16][16] ) );
  DFFRX1 \register_reg[16][15]  ( .D(n1572), .CK(clk), .RN(n2247), .Q(
        \register[16][15] ) );
  DFFRX1 \register_reg[16][14]  ( .D(n1573), .CK(clk), .RN(n2247), .Q(
        \register[16][14] ) );
  DFFRX1 \register_reg[16][13]  ( .D(n1574), .CK(clk), .RN(n2246), .Q(
        \register[16][13] ) );
  DFFRX1 \register_reg[16][12]  ( .D(n1575), .CK(clk), .RN(n2246), .Q(
        \register[16][12] ) );
  DFFRX1 \register_reg[16][11]  ( .D(n1576), .CK(clk), .RN(n2246), .Q(
        \register[16][11] ) );
  DFFRX1 \register_reg[16][10]  ( .D(n1577), .CK(clk), .RN(n2246), .Q(
        \register[16][10] ) );
  DFFRX1 \register_reg[16][9]  ( .D(n1578), .CK(clk), .RN(n2246), .Q(
        \register[16][9] ) );
  DFFRX1 \register_reg[20][31]  ( .D(n1684), .CK(clk), .RN(n2238), .Q(
        \register[20][31] ) );
  DFFRX1 \register_reg[20][30]  ( .D(n1685), .CK(clk), .RN(n2238), .Q(
        \register[20][30] ) );
  DFFRX1 \register_reg[20][29]  ( .D(n1686), .CK(clk), .RN(n2238), .Q(
        \register[20][29] ) );
  DFFRX1 \register_reg[20][28]  ( .D(n1687), .CK(clk), .RN(n2238), .Q(
        \register[20][28] ) );
  DFFRX1 \register_reg[20][27]  ( .D(n1688), .CK(clk), .RN(n2238), .Q(
        \register[20][27] ) );
  DFFRX1 \register_reg[20][26]  ( .D(n1689), .CK(clk), .RN(n2238), .Q(
        \register[20][26] ) );
  DFFRX1 \register_reg[20][25]  ( .D(n1690), .CK(clk), .RN(n2238), .Q(
        \register[20][25] ) );
  DFFRX1 \register_reg[20][24]  ( .D(n1691), .CK(clk), .RN(n2237), .Q(
        \register[20][24] ) );
  DFFRX1 \register_reg[20][23]  ( .D(n1692), .CK(clk), .RN(n2237), .Q(
        \register[20][23] ) );
  DFFRX1 \register_reg[20][22]  ( .D(n1693), .CK(clk), .RN(n2237), .Q(
        \register[20][22] ) );
  DFFRX1 \register_reg[20][21]  ( .D(n1694), .CK(clk), .RN(n2237), .Q(
        \register[20][21] ) );
  DFFRX1 \register_reg[20][20]  ( .D(n1695), .CK(clk), .RN(n2237), .Q(
        \register[20][20] ) );
  DFFRX1 \register_reg[20][19]  ( .D(n1696), .CK(clk), .RN(n2237), .Q(
        \register[20][19] ) );
  DFFRX1 \register_reg[20][18]  ( .D(n1697), .CK(clk), .RN(n2237), .Q(
        \register[20][18] ) );
  DFFRX1 \register_reg[20][17]  ( .D(n1698), .CK(clk), .RN(n2237), .Q(
        \register[20][17] ) );
  DFFRX1 \register_reg[20][16]  ( .D(n1699), .CK(clk), .RN(n2237), .Q(
        \register[20][16] ) );
  DFFRX1 \register_reg[20][15]  ( .D(n1700), .CK(clk), .RN(n2237), .Q(
        \register[20][15] ) );
  DFFRX1 \register_reg[20][14]  ( .D(n1701), .CK(clk), .RN(n2237), .Q(
        \register[20][14] ) );
  DFFRX1 \register_reg[20][13]  ( .D(n1702), .CK(clk), .RN(n2237), .Q(
        \register[20][13] ) );
  DFFRX1 \register_reg[20][12]  ( .D(n1703), .CK(clk), .RN(n2237), .Q(
        \register[20][12] ) );
  DFFRX1 \register_reg[20][11]  ( .D(n1704), .CK(clk), .RN(n2236), .Q(
        \register[20][11] ) );
  DFFRX1 \register_reg[20][10]  ( .D(n1705), .CK(clk), .RN(n2236), .Q(
        \register[20][10] ) );
  DFFRX1 \register_reg[20][9]  ( .D(n1706), .CK(clk), .RN(n2236), .Q(
        \register[20][9] ) );
  DFFRX1 \register_reg[24][31]  ( .D(n1812), .CK(clk), .RN(n2228), .Q(
        \register[24][31] ) );
  DFFRX1 \register_reg[24][30]  ( .D(n1813), .CK(clk), .RN(n2228), .Q(
        \register[24][30] ) );
  DFFRX1 \register_reg[24][29]  ( .D(n1814), .CK(clk), .RN(n2228), .Q(
        \register[24][29] ) );
  DFFRX1 \register_reg[24][28]  ( .D(n1815), .CK(clk), .RN(n2228), .Q(
        \register[24][28] ) );
  DFFRX1 \register_reg[24][27]  ( .D(n1816), .CK(clk), .RN(n2228), .Q(
        \register[24][27] ) );
  DFFRX1 \register_reg[24][26]  ( .D(n1817), .CK(clk), .RN(n2228), .Q(
        \register[24][26] ) );
  DFFRX1 \register_reg[24][25]  ( .D(n1818), .CK(clk), .RN(n2228), .Q(
        \register[24][25] ) );
  DFFRX1 \register_reg[24][24]  ( .D(n1819), .CK(clk), .RN(n2228), .Q(
        \register[24][24] ) );
  DFFRX1 \register_reg[24][23]  ( .D(n1820), .CK(clk), .RN(n2228), .Q(
        \register[24][23] ) );
  DFFRX1 \register_reg[24][22]  ( .D(n1821), .CK(clk), .RN(n2227), .Q(
        \register[24][22] ) );
  DFFRX1 \register_reg[24][21]  ( .D(n1822), .CK(clk), .RN(n2227), .Q(
        \register[24][21] ) );
  DFFRX1 \register_reg[24][20]  ( .D(n1823), .CK(clk), .RN(n2227), .Q(
        \register[24][20] ) );
  DFFRX1 \register_reg[24][19]  ( .D(n1824), .CK(clk), .RN(n2227), .Q(
        \register[24][19] ) );
  DFFRX1 \register_reg[24][18]  ( .D(n1825), .CK(clk), .RN(n2227), .Q(
        \register[24][18] ) );
  DFFRX1 \register_reg[24][17]  ( .D(n1826), .CK(clk), .RN(n2227), .Q(
        \register[24][17] ) );
  DFFRX1 \register_reg[24][16]  ( .D(n1827), .CK(clk), .RN(n2227), .Q(
        \register[24][16] ) );
  DFFRX1 \register_reg[24][15]  ( .D(n1828), .CK(clk), .RN(n2227), .Q(
        \register[24][15] ) );
  DFFRX1 \register_reg[24][14]  ( .D(n1829), .CK(clk), .RN(n2227), .Q(
        \register[24][14] ) );
  DFFRX1 \register_reg[24][13]  ( .D(n1830), .CK(clk), .RN(n2227), .Q(
        \register[24][13] ) );
  DFFRX1 \register_reg[24][12]  ( .D(n1831), .CK(clk), .RN(n2227), .Q(
        \register[24][12] ) );
  DFFRX1 \register_reg[24][11]  ( .D(n1832), .CK(clk), .RN(n2227), .Q(
        \register[24][11] ) );
  DFFRX1 \register_reg[24][10]  ( .D(n1833), .CK(clk), .RN(n2227), .Q(
        \register[24][10] ) );
  DFFRX1 \register_reg[24][9]  ( .D(n1834), .CK(clk), .RN(n2226), .Q(
        \register[24][9] ) );
  DFFRX1 \register_reg[28][31]  ( .D(n1940), .CK(clk), .RN(n2218), .Q(
        \register[28][31] ) );
  DFFRX1 \register_reg[28][30]  ( .D(n1941), .CK(clk), .RN(n2218), .Q(
        \register[28][30] ) );
  DFFRX1 \register_reg[28][29]  ( .D(n1942), .CK(clk), .RN(n2218), .Q(
        \register[28][29] ) );
  DFFRX1 \register_reg[28][28]  ( .D(n1943), .CK(clk), .RN(n2218), .Q(
        \register[28][28] ) );
  DFFRX1 \register_reg[28][27]  ( .D(n1944), .CK(clk), .RN(n2218), .Q(
        \register[28][27] ) );
  DFFRX1 \register_reg[28][26]  ( .D(n1945), .CK(clk), .RN(n2218), .Q(
        \register[28][26] ) );
  DFFRX1 \register_reg[28][25]  ( .D(n1946), .CK(clk), .RN(n2218), .Q(
        \register[28][25] ) );
  DFFRX1 \register_reg[28][24]  ( .D(n1947), .CK(clk), .RN(n2218), .Q(
        \register[28][24] ) );
  DFFRX1 \register_reg[28][23]  ( .D(n1948), .CK(clk), .RN(n2218), .Q(
        \register[28][23] ) );
  DFFRX1 \register_reg[28][22]  ( .D(n1949), .CK(clk), .RN(n2218), .Q(
        \register[28][22] ) );
  DFFRX1 \register_reg[28][21]  ( .D(n1950), .CK(clk), .RN(n2218), .Q(
        \register[28][21] ) );
  DFFRX1 \register_reg[28][20]  ( .D(n1951), .CK(clk), .RN(n2217), .Q(
        \register[28][20] ) );
  DFFRX1 \register_reg[28][19]  ( .D(n1952), .CK(clk), .RN(n2217), .Q(
        \register[28][19] ) );
  DFFRX1 \register_reg[28][18]  ( .D(n1953), .CK(clk), .RN(n2217), .Q(
        \register[28][18] ) );
  DFFRX1 \register_reg[28][17]  ( .D(n1954), .CK(clk), .RN(n2217), .Q(
        \register[28][17] ) );
  DFFRX1 \register_reg[28][16]  ( .D(n1955), .CK(clk), .RN(n2217), .Q(
        \register[28][16] ) );
  DFFRX1 \register_reg[28][15]  ( .D(n1956), .CK(clk), .RN(n2217), .Q(
        \register[28][15] ) );
  DFFRX1 \register_reg[28][14]  ( .D(n1957), .CK(clk), .RN(n2217), .Q(
        \register[28][14] ) );
  DFFRX1 \register_reg[28][13]  ( .D(n1958), .CK(clk), .RN(n2217), .Q(
        \register[28][13] ) );
  DFFRX1 \register_reg[28][12]  ( .D(n1959), .CK(clk), .RN(n2217), .Q(
        \register[28][12] ) );
  DFFRX1 \register_reg[28][11]  ( .D(n1960), .CK(clk), .RN(n2217), .Q(
        \register[28][11] ) );
  DFFRX1 \register_reg[28][10]  ( .D(n1961), .CK(clk), .RN(n2217), .Q(
        \register[28][10] ) );
  DFFRX1 \register_reg[28][9]  ( .D(n1962), .CK(clk), .RN(n2217), .Q(
        \register[28][9] ) );
  DFFRX1 \register_reg[2][31]  ( .D(n1108), .CK(clk), .RN(n2282), .Q(
        \register[2][31] ) );
  DFFRX1 \register_reg[2][30]  ( .D(n1109), .CK(clk), .RN(n2282), .Q(
        \register[2][30] ) );
  DFFRX1 \register_reg[2][29]  ( .D(n1110), .CK(clk), .RN(n2282), .Q(
        \register[2][29] ) );
  DFFRX1 \register_reg[2][28]  ( .D(n1111), .CK(clk), .RN(n2282), .Q(
        \register[2][28] ) );
  DFFRX1 \register_reg[2][27]  ( .D(n1112), .CK(clk), .RN(n2282), .Q(
        \register[2][27] ) );
  DFFRX1 \register_reg[2][26]  ( .D(n1113), .CK(clk), .RN(n2282), .Q(
        \register[2][26] ) );
  DFFRX1 \register_reg[2][25]  ( .D(n1114), .CK(clk), .RN(n2282), .Q(
        \register[2][25] ) );
  DFFRX1 \register_reg[2][24]  ( .D(n1115), .CK(clk), .RN(n2282), .Q(
        \register[2][24] ) );
  DFFRX1 \register_reg[2][23]  ( .D(n1116), .CK(clk), .RN(n2282), .Q(
        \register[2][23] ) );
  DFFRX1 \register_reg[2][22]  ( .D(n1117), .CK(clk), .RN(n2282), .Q(
        \register[2][22] ) );
  DFFRX1 \register_reg[2][21]  ( .D(n1118), .CK(clk), .RN(n2282), .Q(
        \register[2][21] ) );
  DFFRX1 \register_reg[2][20]  ( .D(n1119), .CK(clk), .RN(n2281), .Q(
        \register[2][20] ) );
  DFFRX1 \register_reg[2][19]  ( .D(n1120), .CK(clk), .RN(n2281), .Q(
        \register[2][19] ) );
  DFFRX1 \register_reg[2][18]  ( .D(n1121), .CK(clk), .RN(n2281), .Q(
        \register[2][18] ) );
  DFFRX1 \register_reg[2][17]  ( .D(n1122), .CK(clk), .RN(n2281), .Q(
        \register[2][17] ) );
  DFFRX1 \register_reg[2][16]  ( .D(n1123), .CK(clk), .RN(n2281), .Q(
        \register[2][16] ) );
  DFFRX1 \register_reg[2][15]  ( .D(n1124), .CK(clk), .RN(n2281), .Q(
        \register[2][15] ) );
  DFFRX1 \register_reg[2][14]  ( .D(n1125), .CK(clk), .RN(n2281), .Q(
        \register[2][14] ) );
  DFFRX1 \register_reg[2][13]  ( .D(n1126), .CK(clk), .RN(n2281), .Q(
        \register[2][13] ) );
  DFFRX1 \register_reg[2][12]  ( .D(n1127), .CK(clk), .RN(n2281), .Q(
        \register[2][12] ) );
  DFFRX1 \register_reg[2][11]  ( .D(n1128), .CK(clk), .RN(n2281), .Q(
        \register[2][11] ) );
  DFFRX1 \register_reg[2][10]  ( .D(n1129), .CK(clk), .RN(n2281), .Q(
        \register[2][10] ) );
  DFFRX1 \register_reg[2][9]  ( .D(n1130), .CK(clk), .RN(n2281), .Q(
        \register[2][9] ) );
  DFFRX1 \register_reg[6][31]  ( .D(n1236), .CK(clk), .RN(n2272), .Q(
        \register[6][31] ) );
  DFFRX1 \register_reg[6][30]  ( .D(n1237), .CK(clk), .RN(n2272), .Q(
        \register[6][30] ) );
  DFFRX1 \register_reg[6][29]  ( .D(n1238), .CK(clk), .RN(n2272), .Q(
        \register[6][29] ) );
  DFFRX1 \register_reg[6][28]  ( .D(n1239), .CK(clk), .RN(n2272), .Q(
        \register[6][28] ) );
  DFFRX1 \register_reg[6][27]  ( .D(n1240), .CK(clk), .RN(n2272), .Q(
        \register[6][27] ) );
  DFFRX1 \register_reg[6][26]  ( .D(n1241), .CK(clk), .RN(n2272), .Q(
        \register[6][26] ) );
  DFFRX1 \register_reg[6][25]  ( .D(n1242), .CK(clk), .RN(n2272), .Q(
        \register[6][25] ) );
  DFFRX1 \register_reg[6][24]  ( .D(n1243), .CK(clk), .RN(n2272), .Q(
        \register[6][24] ) );
  DFFRX1 \register_reg[6][23]  ( .D(n1244), .CK(clk), .RN(n2272), .Q(
        \register[6][23] ) );
  DFFRX1 \register_reg[6][22]  ( .D(n1245), .CK(clk), .RN(n2272), .Q(
        \register[6][22] ) );
  DFFRX1 \register_reg[6][21]  ( .D(n1246), .CK(clk), .RN(n2272), .Q(
        \register[6][21] ) );
  DFFRX1 \register_reg[6][20]  ( .D(n1247), .CK(clk), .RN(n2272), .Q(
        \register[6][20] ) );
  DFFRX1 \register_reg[6][19]  ( .D(n1248), .CK(clk), .RN(n2272), .Q(
        \register[6][19] ) );
  DFFRX1 \register_reg[6][18]  ( .D(n1249), .CK(clk), .RN(n2271), .Q(
        \register[6][18] ) );
  DFFRX1 \register_reg[6][17]  ( .D(n1250), .CK(clk), .RN(n2271), .Q(
        \register[6][17] ) );
  DFFRX1 \register_reg[6][16]  ( .D(n1251), .CK(clk), .RN(n2271), .Q(
        \register[6][16] ) );
  DFFRX1 \register_reg[6][15]  ( .D(n1252), .CK(clk), .RN(n2271), .Q(
        \register[6][15] ) );
  DFFRX1 \register_reg[6][14]  ( .D(n1253), .CK(clk), .RN(n2271), .Q(
        \register[6][14] ) );
  DFFRX1 \register_reg[6][13]  ( .D(n1254), .CK(clk), .RN(n2271), .Q(
        \register[6][13] ) );
  DFFRX1 \register_reg[6][12]  ( .D(n1255), .CK(clk), .RN(n2271), .Q(
        \register[6][12] ) );
  DFFRX1 \register_reg[6][11]  ( .D(n1256), .CK(clk), .RN(n2271), .Q(
        \register[6][11] ) );
  DFFRX1 \register_reg[6][10]  ( .D(n1257), .CK(clk), .RN(n2271), .Q(
        \register[6][10] ) );
  DFFRX1 \register_reg[6][9]  ( .D(n1258), .CK(clk), .RN(n2271), .Q(
        \register[6][9] ) );
  DFFRX1 \register_reg[10][31]  ( .D(n1364), .CK(clk), .RN(n2263), .Q(
        \register[10][31] ) );
  DFFRX1 \register_reg[10][30]  ( .D(n1365), .CK(clk), .RN(n2263), .Q(
        \register[10][30] ) );
  DFFRX1 \register_reg[10][29]  ( .D(n1366), .CK(clk), .RN(n2262), .Q(
        \register[10][29] ) );
  DFFRX1 \register_reg[10][28]  ( .D(n1367), .CK(clk), .RN(n2262), .Q(
        \register[10][28] ) );
  DFFRX1 \register_reg[10][27]  ( .D(n1368), .CK(clk), .RN(n2262), .Q(
        \register[10][27] ) );
  DFFRX1 \register_reg[10][26]  ( .D(n1369), .CK(clk), .RN(n2262), .Q(
        \register[10][26] ) );
  DFFRX1 \register_reg[10][25]  ( .D(n1370), .CK(clk), .RN(n2262), .Q(
        \register[10][25] ) );
  DFFRX1 \register_reg[10][24]  ( .D(n1371), .CK(clk), .RN(n2262), .Q(
        \register[10][24] ) );
  DFFRX1 \register_reg[10][23]  ( .D(n1372), .CK(clk), .RN(n2262), .Q(
        \register[10][23] ) );
  DFFRX1 \register_reg[10][22]  ( .D(n1373), .CK(clk), .RN(n2262), .Q(
        \register[10][22] ) );
  DFFRX1 \register_reg[10][21]  ( .D(n1374), .CK(clk), .RN(n2262), .Q(
        \register[10][21] ) );
  DFFRX1 \register_reg[10][20]  ( .D(n1375), .CK(clk), .RN(n2262), .Q(
        \register[10][20] ) );
  DFFRX1 \register_reg[10][19]  ( .D(n1376), .CK(clk), .RN(n2262), .Q(
        \register[10][19] ) );
  DFFRX1 \register_reg[10][18]  ( .D(n1377), .CK(clk), .RN(n2262), .Q(
        \register[10][18] ) );
  DFFRX1 \register_reg[10][17]  ( .D(n1378), .CK(clk), .RN(n2262), .Q(
        \register[10][17] ) );
  DFFRX1 \register_reg[10][16]  ( .D(n1379), .CK(clk), .RN(n2261), .Q(
        \register[10][16] ) );
  DFFRX1 \register_reg[10][15]  ( .D(n1380), .CK(clk), .RN(n2261), .Q(
        \register[10][15] ) );
  DFFRX1 \register_reg[10][14]  ( .D(n1381), .CK(clk), .RN(n2261), .Q(
        \register[10][14] ) );
  DFFRX1 \register_reg[10][13]  ( .D(n1382), .CK(clk), .RN(n2261), .Q(
        \register[10][13] ) );
  DFFRX1 \register_reg[10][12]  ( .D(n1383), .CK(clk), .RN(n2261), .Q(
        \register[10][12] ) );
  DFFRX1 \register_reg[10][11]  ( .D(n1384), .CK(clk), .RN(n2261), .Q(
        \register[10][11] ) );
  DFFRX1 \register_reg[10][10]  ( .D(n1385), .CK(clk), .RN(n2261), .Q(
        \register[10][10] ) );
  DFFRX1 \register_reg[10][9]  ( .D(n1386), .CK(clk), .RN(n2261), .Q(
        \register[10][9] ) );
  DFFRX1 \register_reg[14][31]  ( .D(n1492), .CK(clk), .RN(n2253), .Q(
        \register[14][31] ) );
  DFFRX1 \register_reg[14][30]  ( .D(n1493), .CK(clk), .RN(n2253), .Q(
        \register[14][30] ) );
  DFFRX1 \register_reg[14][29]  ( .D(n1494), .CK(clk), .RN(n2253), .Q(
        \register[14][29] ) );
  DFFRX1 \register_reg[14][28]  ( .D(n1495), .CK(clk), .RN(n2253), .Q(
        \register[14][28] ) );
  DFFRX1 \register_reg[14][27]  ( .D(n1496), .CK(clk), .RN(n2252), .Q(
        \register[14][27] ) );
  DFFRX1 \register_reg[14][26]  ( .D(n1497), .CK(clk), .RN(n2252), .Q(
        \register[14][26] ) );
  DFFRX1 \register_reg[14][25]  ( .D(n1498), .CK(clk), .RN(n2252), .Q(
        \register[14][25] ) );
  DFFRX1 \register_reg[14][24]  ( .D(n1499), .CK(clk), .RN(n2252), .Q(
        \register[14][24] ) );
  DFFRX1 \register_reg[14][23]  ( .D(n1500), .CK(clk), .RN(n2252), .Q(
        \register[14][23] ) );
  DFFRX1 \register_reg[14][22]  ( .D(n1501), .CK(clk), .RN(n2252), .Q(
        \register[14][22] ) );
  DFFRX1 \register_reg[14][21]  ( .D(n1502), .CK(clk), .RN(n2252), .Q(
        \register[14][21] ) );
  DFFRX1 \register_reg[14][20]  ( .D(n1503), .CK(clk), .RN(n2252), .Q(
        \register[14][20] ) );
  DFFRX1 \register_reg[14][19]  ( .D(n1504), .CK(clk), .RN(n2252), .Q(
        \register[14][19] ) );
  DFFRX1 \register_reg[14][18]  ( .D(n1505), .CK(clk), .RN(n2252), .Q(
        \register[14][18] ) );
  DFFRX1 \register_reg[14][17]  ( .D(n1506), .CK(clk), .RN(n2252), .Q(
        \register[14][17] ) );
  DFFRX1 \register_reg[14][16]  ( .D(n1507), .CK(clk), .RN(n2252), .Q(
        \register[14][16] ) );
  DFFRX1 \register_reg[14][15]  ( .D(n1508), .CK(clk), .RN(n2252), .Q(
        \register[14][15] ) );
  DFFRX1 \register_reg[14][14]  ( .D(n1509), .CK(clk), .RN(n2251), .Q(
        \register[14][14] ) );
  DFFRX1 \register_reg[14][13]  ( .D(n1510), .CK(clk), .RN(n2251), .Q(
        \register[14][13] ) );
  DFFRX1 \register_reg[14][12]  ( .D(n1511), .CK(clk), .RN(n2251), .Q(
        \register[14][12] ) );
  DFFRX1 \register_reg[14][11]  ( .D(n1512), .CK(clk), .RN(n2251), .Q(
        \register[14][11] ) );
  DFFRX1 \register_reg[14][10]  ( .D(n1513), .CK(clk), .RN(n2251), .Q(
        \register[14][10] ) );
  DFFRX1 \register_reg[14][9]  ( .D(n1514), .CK(clk), .RN(n2251), .Q(
        \register[14][9] ) );
  DFFRX1 \register_reg[18][31]  ( .D(n1620), .CK(clk), .RN(n2243), .Q(
        \register[18][31] ) );
  DFFRX1 \register_reg[18][30]  ( .D(n1621), .CK(clk), .RN(n2243), .Q(
        \register[18][30] ) );
  DFFRX1 \register_reg[18][29]  ( .D(n1622), .CK(clk), .RN(n2243), .Q(
        \register[18][29] ) );
  DFFRX1 \register_reg[18][28]  ( .D(n1623), .CK(clk), .RN(n2243), .Q(
        \register[18][28] ) );
  DFFRX1 \register_reg[18][27]  ( .D(n1624), .CK(clk), .RN(n2243), .Q(
        \register[18][27] ) );
  DFFRX1 \register_reg[18][26]  ( .D(n1625), .CK(clk), .RN(n2243), .Q(
        \register[18][26] ) );
  DFFRX1 \register_reg[18][25]  ( .D(n1626), .CK(clk), .RN(n2242), .Q(
        \register[18][25] ) );
  DFFRX1 \register_reg[18][24]  ( .D(n1627), .CK(clk), .RN(n2242), .Q(
        \register[18][24] ) );
  DFFRX1 \register_reg[18][23]  ( .D(n1628), .CK(clk), .RN(n2242), .Q(
        \register[18][23] ) );
  DFFRX1 \register_reg[18][22]  ( .D(n1629), .CK(clk), .RN(n2242), .Q(
        \register[18][22] ) );
  DFFRX1 \register_reg[18][21]  ( .D(n1630), .CK(clk), .RN(n2242), .Q(
        \register[18][21] ) );
  DFFRX1 \register_reg[18][20]  ( .D(n1631), .CK(clk), .RN(n2242), .Q(
        \register[18][20] ) );
  DFFRX1 \register_reg[18][19]  ( .D(n1632), .CK(clk), .RN(n2242), .Q(
        \register[18][19] ) );
  DFFRX1 \register_reg[18][18]  ( .D(n1633), .CK(clk), .RN(n2242), .Q(
        \register[18][18] ) );
  DFFRX1 \register_reg[18][17]  ( .D(n1634), .CK(clk), .RN(n2242), .Q(
        \register[18][17] ) );
  DFFRX1 \register_reg[18][16]  ( .D(n1635), .CK(clk), .RN(n2242), .Q(
        \register[18][16] ) );
  DFFRX1 \register_reg[18][15]  ( .D(n1636), .CK(clk), .RN(n2242), .Q(
        \register[18][15] ) );
  DFFRX1 \register_reg[18][14]  ( .D(n1637), .CK(clk), .RN(n2242), .Q(
        \register[18][14] ) );
  DFFRX1 \register_reg[18][13]  ( .D(n1638), .CK(clk), .RN(n2242), .Q(
        \register[18][13] ) );
  DFFRX1 \register_reg[18][12]  ( .D(n1639), .CK(clk), .RN(n2241), .Q(
        \register[18][12] ) );
  DFFRX1 \register_reg[18][11]  ( .D(n1640), .CK(clk), .RN(n2241), .Q(
        \register[18][11] ) );
  DFFRX1 \register_reg[18][10]  ( .D(n1641), .CK(clk), .RN(n2241), .Q(
        \register[18][10] ) );
  DFFRX1 \register_reg[18][9]  ( .D(n1642), .CK(clk), .RN(n2241), .Q(
        \register[18][9] ) );
  DFFRX1 \register_reg[22][31]  ( .D(n1748), .CK(clk), .RN(n2233), .Q(
        \register[22][31] ) );
  DFFRX1 \register_reg[22][30]  ( .D(n1749), .CK(clk), .RN(n2233), .Q(
        \register[22][30] ) );
  DFFRX1 \register_reg[22][29]  ( .D(n1750), .CK(clk), .RN(n2233), .Q(
        \register[22][29] ) );
  DFFRX1 \register_reg[22][28]  ( .D(n1751), .CK(clk), .RN(n2233), .Q(
        \register[22][28] ) );
  DFFRX1 \register_reg[22][27]  ( .D(n1752), .CK(clk), .RN(n2233), .Q(
        \register[22][27] ) );
  DFFRX1 \register_reg[22][26]  ( .D(n1753), .CK(clk), .RN(n2233), .Q(
        \register[22][26] ) );
  DFFRX1 \register_reg[22][25]  ( .D(n1754), .CK(clk), .RN(n2233), .Q(
        \register[22][25] ) );
  DFFRX1 \register_reg[22][24]  ( .D(n1755), .CK(clk), .RN(n2233), .Q(
        \register[22][24] ) );
  DFFRX1 \register_reg[22][23]  ( .D(n1756), .CK(clk), .RN(n2232), .Q(
        \register[22][23] ) );
  DFFRX1 \register_reg[22][22]  ( .D(n1757), .CK(clk), .RN(n2232), .Q(
        \register[22][22] ) );
  DFFRX1 \register_reg[22][21]  ( .D(n1758), .CK(clk), .RN(n2232), .Q(
        \register[22][21] ) );
  DFFRX1 \register_reg[22][20]  ( .D(n1759), .CK(clk), .RN(n2232), .Q(
        \register[22][20] ) );
  DFFRX1 \register_reg[22][19]  ( .D(n1760), .CK(clk), .RN(n2232), .Q(
        \register[22][19] ) );
  DFFRX1 \register_reg[22][18]  ( .D(n1761), .CK(clk), .RN(n2232), .Q(
        \register[22][18] ) );
  DFFRX1 \register_reg[22][17]  ( .D(n1762), .CK(clk), .RN(n2232), .Q(
        \register[22][17] ) );
  DFFRX1 \register_reg[22][16]  ( .D(n1763), .CK(clk), .RN(n2232), .Q(
        \register[22][16] ) );
  DFFRX1 \register_reg[22][15]  ( .D(n1764), .CK(clk), .RN(n2232), .Q(
        \register[22][15] ) );
  DFFRX1 \register_reg[22][14]  ( .D(n1765), .CK(clk), .RN(n2232), .Q(
        \register[22][14] ) );
  DFFRX1 \register_reg[22][13]  ( .D(n1766), .CK(clk), .RN(n2232), .Q(
        \register[22][13] ) );
  DFFRX1 \register_reg[22][12]  ( .D(n1767), .CK(clk), .RN(n2232), .Q(
        \register[22][12] ) );
  DFFRX1 \register_reg[22][11]  ( .D(n1768), .CK(clk), .RN(n2232), .Q(
        \register[22][11] ) );
  DFFRX1 \register_reg[22][10]  ( .D(n1769), .CK(clk), .RN(n2231), .Q(
        \register[22][10] ) );
  DFFRX1 \register_reg[22][9]  ( .D(n1770), .CK(clk), .RN(n2231), .Q(
        \register[22][9] ) );
  DFFRX1 \register_reg[26][31]  ( .D(n1876), .CK(clk), .RN(n2223), .Q(
        \register[26][31] ) );
  DFFRX1 \register_reg[26][30]  ( .D(n1877), .CK(clk), .RN(n2223), .Q(
        \register[26][30] ) );
  DFFRX1 \register_reg[26][29]  ( .D(n1878), .CK(clk), .RN(n2223), .Q(
        \register[26][29] ) );
  DFFRX1 \register_reg[26][28]  ( .D(n1879), .CK(clk), .RN(n2223), .Q(
        \register[26][28] ) );
  DFFRX1 \register_reg[26][27]  ( .D(n1880), .CK(clk), .RN(n2223), .Q(
        \register[26][27] ) );
  DFFRX1 \register_reg[26][26]  ( .D(n1881), .CK(clk), .RN(n2223), .Q(
        \register[26][26] ) );
  DFFRX1 \register_reg[26][25]  ( .D(n1882), .CK(clk), .RN(n2223), .Q(
        \register[26][25] ) );
  DFFRX1 \register_reg[26][24]  ( .D(n1883), .CK(clk), .RN(n2223), .Q(
        \register[26][24] ) );
  DFFRX1 \register_reg[26][23]  ( .D(n1884), .CK(clk), .RN(n2223), .Q(
        \register[26][23] ) );
  DFFRX1 \register_reg[26][22]  ( .D(n1885), .CK(clk), .RN(n2223), .Q(
        \register[26][22] ) );
  DFFRX1 \register_reg[26][21]  ( .D(n1886), .CK(clk), .RN(n2222), .Q(
        \register[26][21] ) );
  DFFRX1 \register_reg[26][20]  ( .D(n1887), .CK(clk), .RN(n2222), .Q(
        \register[26][20] ) );
  DFFRX1 \register_reg[26][19]  ( .D(n1888), .CK(clk), .RN(n2222), .Q(
        \register[26][19] ) );
  DFFRX1 \register_reg[26][18]  ( .D(n1889), .CK(clk), .RN(n2222), .Q(
        \register[26][18] ) );
  DFFRX1 \register_reg[26][17]  ( .D(n1890), .CK(clk), .RN(n2222), .Q(
        \register[26][17] ) );
  DFFRX1 \register_reg[26][16]  ( .D(n1891), .CK(clk), .RN(n2222), .Q(
        \register[26][16] ) );
  DFFRX1 \register_reg[26][15]  ( .D(n1892), .CK(clk), .RN(n2222), .Q(
        \register[26][15] ) );
  DFFRX1 \register_reg[26][14]  ( .D(n1893), .CK(clk), .RN(n2222), .Q(
        \register[26][14] ) );
  DFFRX1 \register_reg[26][13]  ( .D(n1894), .CK(clk), .RN(n2222), .Q(
        \register[26][13] ) );
  DFFRX1 \register_reg[26][12]  ( .D(n1895), .CK(clk), .RN(n2222), .Q(
        \register[26][12] ) );
  DFFRX1 \register_reg[26][11]  ( .D(n1896), .CK(clk), .RN(n2222), .Q(
        \register[26][11] ) );
  DFFRX1 \register_reg[26][10]  ( .D(n1897), .CK(clk), .RN(n2222), .Q(
        \register[26][10] ) );
  DFFRX1 \register_reg[26][9]  ( .D(n1898), .CK(clk), .RN(n2222), .Q(
        \register[26][9] ) );
  DFFRX1 \register_reg[30][31]  ( .D(n2004), .CK(clk), .RN(n2213), .Q(
        \register[30][31] ) );
  DFFRX1 \register_reg[30][30]  ( .D(n2005), .CK(clk), .RN(n2213), .Q(
        \register[30][30] ) );
  DFFRX1 \register_reg[30][29]  ( .D(n2006), .CK(clk), .RN(n2213), .Q(
        \register[30][29] ) );
  DFFRX1 \register_reg[30][28]  ( .D(n2007), .CK(clk), .RN(n2213), .Q(
        \register[30][28] ) );
  DFFRX1 \register_reg[30][27]  ( .D(n2008), .CK(clk), .RN(n2213), .Q(
        \register[30][27] ) );
  DFFRX1 \register_reg[30][26]  ( .D(n2009), .CK(clk), .RN(n2213), .Q(
        \register[30][26] ) );
  DFFRX1 \register_reg[30][25]  ( .D(n2010), .CK(clk), .RN(n2213), .Q(
        \register[30][25] ) );
  DFFRX1 \register_reg[30][24]  ( .D(n2011), .CK(clk), .RN(n2213), .Q(
        \register[30][24] ) );
  DFFRX1 \register_reg[30][23]  ( .D(n2012), .CK(clk), .RN(n2213), .Q(
        \register[30][23] ) );
  DFFRX1 \register_reg[30][22]  ( .D(n2013), .CK(clk), .RN(n2213), .Q(
        \register[30][22] ) );
  DFFRX1 \register_reg[30][21]  ( .D(n2014), .CK(clk), .RN(n2213), .Q(
        \register[30][21] ) );
  DFFRX1 \register_reg[30][20]  ( .D(n2015), .CK(clk), .RN(n2213), .Q(
        \register[30][20] ) );
  DFFRX1 \register_reg[30][19]  ( .D(n2016), .CK(clk), .RN(n2212), .Q(
        \register[30][19] ) );
  DFFRX1 \register_reg[30][18]  ( .D(n2017), .CK(clk), .RN(n2212), .Q(
        \register[30][18] ) );
  DFFRX1 \register_reg[30][17]  ( .D(n2018), .CK(clk), .RN(n2212), .Q(
        \register[30][17] ) );
  DFFRX1 \register_reg[30][16]  ( .D(n2019), .CK(clk), .RN(n2212), .Q(
        \register[30][16] ) );
  DFFRX1 \register_reg[30][15]  ( .D(n2020), .CK(clk), .RN(n2212), .Q(
        \register[30][15] ) );
  DFFRX1 \register_reg[30][14]  ( .D(n2021), .CK(clk), .RN(n2212), .Q(
        \register[30][14] ) );
  DFFRX1 \register_reg[30][13]  ( .D(n2022), .CK(clk), .RN(n2212), .Q(
        \register[30][13] ) );
  DFFRX1 \register_reg[30][12]  ( .D(n2023), .CK(clk), .RN(n2212), .Q(
        \register[30][12] ) );
  DFFRX1 \register_reg[30][11]  ( .D(n2024), .CK(clk), .RN(n2212), .Q(
        \register[30][11] ) );
  DFFRX1 \register_reg[30][10]  ( .D(n2025), .CK(clk), .RN(n2212), .Q(
        \register[30][10] ) );
  DFFRX1 \register_reg[30][9]  ( .D(n2026), .CK(clk), .RN(n2212), .Q(
        \register[30][9] ) );
  DFFRX1 \register_reg[3][8]  ( .D(n1163), .CK(clk), .RN(n2278), .Q(
        \register[3][8] ) );
  DFFRX1 \register_reg[3][7]  ( .D(n1164), .CK(clk), .RN(n2278), .Q(
        \register[3][7] ) );
  DFFRX1 \register_reg[3][6]  ( .D(n1165), .CK(clk), .RN(n2278), .Q(
        \register[3][6] ) );
  DFFRX1 \register_reg[3][5]  ( .D(n1166), .CK(clk), .RN(n2278), .Q(
        \register[3][5] ) );
  DFFRX1 \register_reg[3][4]  ( .D(n1167), .CK(clk), .RN(n2278), .Q(
        \register[3][4] ) );
  DFFRX1 \register_reg[7][8]  ( .D(n1291), .CK(clk), .RN(n2268), .Q(
        \register[7][8] ) );
  DFFRX1 \register_reg[7][7]  ( .D(n1292), .CK(clk), .RN(n2268), .Q(
        \register[7][7] ) );
  DFFRX1 \register_reg[7][6]  ( .D(n1293), .CK(clk), .RN(n2268), .Q(
        \register[7][6] ) );
  DFFRX1 \register_reg[7][5]  ( .D(n1294), .CK(clk), .RN(n2268), .Q(
        \register[7][5] ) );
  DFFRX1 \register_reg[7][4]  ( .D(n1295), .CK(clk), .RN(n2268), .Q(
        \register[7][4] ) );
  DFFRX1 \register_reg[11][8]  ( .D(n1419), .CK(clk), .RN(n2258), .Q(
        \register[11][8] ) );
  DFFRX1 \register_reg[11][7]  ( .D(n1420), .CK(clk), .RN(n2258), .Q(
        \register[11][7] ) );
  DFFRX1 \register_reg[11][6]  ( .D(n1421), .CK(clk), .RN(n2258), .Q(
        \register[11][6] ) );
  DFFRX1 \register_reg[11][5]  ( .D(n1422), .CK(clk), .RN(n2258), .Q(
        \register[11][5] ) );
  DFFRX1 \register_reg[11][4]  ( .D(n1423), .CK(clk), .RN(n2258), .Q(
        \register[11][4] ) );
  DFFRX1 \register_reg[15][8]  ( .D(n1547), .CK(clk), .RN(n2249), .Q(
        \register[15][8] ) );
  DFFRX1 \register_reg[15][7]  ( .D(n1548), .CK(clk), .RN(n2248), .Q(
        \register[15][7] ) );
  DFFRX1 \register_reg[15][6]  ( .D(n1549), .CK(clk), .RN(n2248), .Q(
        \register[15][6] ) );
  DFFRX1 \register_reg[15][5]  ( .D(n1550), .CK(clk), .RN(n2248), .Q(
        \register[15][5] ) );
  DFFRX1 \register_reg[15][4]  ( .D(n1551), .CK(clk), .RN(n2248), .Q(
        \register[15][4] ) );
  DFFRX1 \register_reg[19][8]  ( .D(n1675), .CK(clk), .RN(n2239), .Q(
        \register[19][8] ) );
  DFFRX1 \register_reg[19][7]  ( .D(n1676), .CK(clk), .RN(n2239), .Q(
        \register[19][7] ) );
  DFFRX1 \register_reg[19][6]  ( .D(n1677), .CK(clk), .RN(n2239), .Q(
        \register[19][6] ) );
  DFFRX1 \register_reg[19][5]  ( .D(n1678), .CK(clk), .RN(n2238), .Q(
        \register[19][5] ) );
  DFFRX1 \register_reg[19][4]  ( .D(n1679), .CK(clk), .RN(n2238), .Q(
        \register[19][4] ) );
  DFFRX1 \register_reg[23][8]  ( .D(n1803), .CK(clk), .RN(n2229), .Q(
        \register[23][8] ) );
  DFFRX1 \register_reg[23][7]  ( .D(n1804), .CK(clk), .RN(n2229), .Q(
        \register[23][7] ) );
  DFFRX1 \register_reg[23][6]  ( .D(n1805), .CK(clk), .RN(n2229), .Q(
        \register[23][6] ) );
  DFFRX1 \register_reg[23][5]  ( .D(n1806), .CK(clk), .RN(n2229), .Q(
        \register[23][5] ) );
  DFFRX1 \register_reg[23][4]  ( .D(n1807), .CK(clk), .RN(n2229), .Q(
        \register[23][4] ) );
  DFFRX1 \register_reg[27][8]  ( .D(n1931), .CK(clk), .RN(n2219), .Q(
        \register[27][8] ) );
  DFFRX1 \register_reg[27][7]  ( .D(n1932), .CK(clk), .RN(n2219), .Q(
        \register[27][7] ) );
  DFFRX1 \register_reg[27][6]  ( .D(n1933), .CK(clk), .RN(n2219), .Q(
        \register[27][6] ) );
  DFFRX1 \register_reg[27][5]  ( .D(n1934), .CK(clk), .RN(n2219), .Q(
        \register[27][5] ) );
  DFFRX1 \register_reg[27][4]  ( .D(n1935), .CK(clk), .RN(n2219), .Q(
        \register[27][4] ) );
  DFFRX1 \register_reg[31][8]  ( .D(n2059), .CK(clk), .RN(n2209), .Q(
        \register[31][8] ) );
  DFFRX1 \register_reg[31][7]  ( .D(n2060), .CK(clk), .RN(n2209), .Q(
        \register[31][7] ) );
  DFFRX1 \register_reg[31][6]  ( .D(n2061), .CK(clk), .RN(n2209), .Q(
        \register[31][6] ) );
  DFFRX1 \register_reg[31][5]  ( .D(n2062), .CK(clk), .RN(n2209), .Q(
        \register[31][5] ) );
  DFFRX1 \register_reg[31][4]  ( .D(n2063), .CK(clk), .RN(n2209), .Q(
        \register[31][4] ) );
  DFFRX1 \register_reg[3][3]  ( .D(n1168), .CK(clk), .RN(n2278), .Q(
        \register[3][3] ) );
  DFFRX1 \register_reg[3][2]  ( .D(n1169), .CK(clk), .RN(n2278), .Q(
        \register[3][2] ) );
  DFFRX1 \register_reg[3][1]  ( .D(n1170), .CK(clk), .RN(n2278), .Q(
        \register[3][1] ) );
  DFFRX1 \register_reg[3][0]  ( .D(n1171), .CK(clk), .RN(n2277), .Q(
        \register[3][0] ) );
  DFFRX1 \register_reg[7][3]  ( .D(n1296), .CK(clk), .RN(n2268), .Q(
        \register[7][3] ) );
  DFFRX1 \register_reg[7][2]  ( .D(n1297), .CK(clk), .RN(n2268), .Q(
        \register[7][2] ) );
  DFFRX1 \register_reg[7][1]  ( .D(n1298), .CK(clk), .RN(n2268), .Q(
        \register[7][1] ) );
  DFFRX1 \register_reg[7][0]  ( .D(n1299), .CK(clk), .RN(n2268), .Q(
        \register[7][0] ) );
  DFFRX1 \register_reg[11][3]  ( .D(n1424), .CK(clk), .RN(n2258), .Q(
        \register[11][3] ) );
  DFFRX1 \register_reg[11][2]  ( .D(n1425), .CK(clk), .RN(n2258), .Q(
        \register[11][2] ) );
  DFFRX1 \register_reg[11][1]  ( .D(n1426), .CK(clk), .RN(n2258), .Q(
        \register[11][1] ) );
  DFFRX1 \register_reg[11][0]  ( .D(n1427), .CK(clk), .RN(n2258), .Q(
        \register[11][0] ) );
  DFFRX1 \register_reg[15][3]  ( .D(n1552), .CK(clk), .RN(n2248), .Q(
        \register[15][3] ) );
  DFFRX1 \register_reg[15][2]  ( .D(n1553), .CK(clk), .RN(n2248), .Q(
        \register[15][2] ) );
  DFFRX1 \register_reg[15][1]  ( .D(n1554), .CK(clk), .RN(n2248), .Q(
        \register[15][1] ) );
  DFFRX1 \register_reg[15][0]  ( .D(n1555), .CK(clk), .RN(n2248), .Q(
        \register[15][0] ) );
  DFFRX1 \register_reg[19][3]  ( .D(n1680), .CK(clk), .RN(n2238), .Q(
        \register[19][3] ) );
  DFFRX1 \register_reg[19][2]  ( .D(n1681), .CK(clk), .RN(n2238), .Q(
        \register[19][2] ) );
  DFFRX1 \register_reg[19][1]  ( .D(n1682), .CK(clk), .RN(n2238), .Q(
        \register[19][1] ) );
  DFFRX1 \register_reg[19][0]  ( .D(n1683), .CK(clk), .RN(n2238), .Q(
        \register[19][0] ) );
  DFFRX1 \register_reg[23][3]  ( .D(n1808), .CK(clk), .RN(n2228), .Q(
        \register[23][3] ) );
  DFFRX1 \register_reg[23][2]  ( .D(n1809), .CK(clk), .RN(n2228), .Q(
        \register[23][2] ) );
  DFFRX1 \register_reg[23][1]  ( .D(n1810), .CK(clk), .RN(n2228), .Q(
        \register[23][1] ) );
  DFFRX1 \register_reg[23][0]  ( .D(n1811), .CK(clk), .RN(n2228), .Q(
        \register[23][0] ) );
  DFFRX1 \register_reg[27][3]  ( .D(n1936), .CK(clk), .RN(n2219), .Q(
        \register[27][3] ) );
  DFFRX1 \register_reg[27][2]  ( .D(n1937), .CK(clk), .RN(n2219), .Q(
        \register[27][2] ) );
  DFFRX1 \register_reg[27][1]  ( .D(n1938), .CK(clk), .RN(n2218), .Q(
        \register[27][1] ) );
  DFFRX1 \register_reg[27][0]  ( .D(n1939), .CK(clk), .RN(n2218), .Q(
        \register[27][0] ) );
  DFFRX1 \register_reg[31][3]  ( .D(n2064), .CK(clk), .RN(n2209), .Q(
        \register[31][3] ) );
  DFFRX1 \register_reg[31][1]  ( .D(n2066), .CK(clk), .RN(n2209), .Q(
        \register[31][1] ) );
  DFFRX1 \register_reg[31][2]  ( .D(n2065), .CK(clk), .RN(n2209), .Q(
        \register[31][2] ) );
  DFFRX1 \register_reg[1][8]  ( .D(n1099), .CK(clk), .RN(n2283), .Q(
        \register[1][8] ) );
  DFFRX1 \register_reg[1][7]  ( .D(n1100), .CK(clk), .RN(n2283), .Q(
        \register[1][7] ) );
  DFFRX1 \register_reg[1][6]  ( .D(n1101), .CK(clk), .RN(n2283), .Q(
        \register[1][6] ) );
  DFFRX1 \register_reg[1][5]  ( .D(n1102), .CK(clk), .RN(n2283), .Q(
        \register[1][5] ) );
  DFFRX1 \register_reg[1][4]  ( .D(n1103), .CK(clk), .RN(n2283), .Q(
        \register[1][4] ) );
  DFFRX1 \register_reg[5][8]  ( .D(n1227), .CK(clk), .RN(n2273), .Q(
        \register[5][8] ) );
  DFFRX1 \register_reg[5][7]  ( .D(n1228), .CK(clk), .RN(n2273), .Q(
        \register[5][7] ) );
  DFFRX1 \register_reg[5][6]  ( .D(n1229), .CK(clk), .RN(n2273), .Q(
        \register[5][6] ) );
  DFFRX1 \register_reg[5][5]  ( .D(n1230), .CK(clk), .RN(n2273), .Q(
        \register[5][5] ) );
  DFFRX1 \register_reg[5][4]  ( .D(n1231), .CK(clk), .RN(n2273), .Q(
        \register[5][4] ) );
  DFFRX1 \register_reg[9][8]  ( .D(n1355), .CK(clk), .RN(n2263), .Q(
        \register[9][8] ) );
  DFFRX1 \register_reg[9][7]  ( .D(n1356), .CK(clk), .RN(n2263), .Q(
        \register[9][7] ) );
  DFFRX1 \register_reg[9][6]  ( .D(n1357), .CK(clk), .RN(n2263), .Q(
        \register[9][6] ) );
  DFFRX1 \register_reg[9][5]  ( .D(n1358), .CK(clk), .RN(n2263), .Q(
        \register[9][5] ) );
  DFFRX1 \register_reg[9][4]  ( .D(n1359), .CK(clk), .RN(n2263), .Q(
        \register[9][4] ) );
  DFFRX1 \register_reg[13][8]  ( .D(n1483), .CK(clk), .RN(n2253), .Q(
        \register[13][8] ) );
  DFFRX1 \register_reg[13][7]  ( .D(n1484), .CK(clk), .RN(n2253), .Q(
        \register[13][7] ) );
  DFFRX1 \register_reg[13][6]  ( .D(n1485), .CK(clk), .RN(n2253), .Q(
        \register[13][6] ) );
  DFFRX1 \register_reg[13][5]  ( .D(n1486), .CK(clk), .RN(n2253), .Q(
        \register[13][5] ) );
  DFFRX1 \register_reg[13][4]  ( .D(n1487), .CK(clk), .RN(n2253), .Q(
        \register[13][4] ) );
  DFFRX1 \register_reg[17][8]  ( .D(n1611), .CK(clk), .RN(n2244), .Q(
        \register[17][8] ) );
  DFFRX1 \register_reg[17][7]  ( .D(n1612), .CK(clk), .RN(n2244), .Q(
        \register[17][7] ) );
  DFFRX1 \register_reg[17][6]  ( .D(n1613), .CK(clk), .RN(n2243), .Q(
        \register[17][6] ) );
  DFFRX1 \register_reg[17][5]  ( .D(n1614), .CK(clk), .RN(n2243), .Q(
        \register[17][5] ) );
  DFFRX1 \register_reg[17][4]  ( .D(n1615), .CK(clk), .RN(n2243), .Q(
        \register[17][4] ) );
  DFFRX1 \register_reg[21][8]  ( .D(n1739), .CK(clk), .RN(n2234), .Q(
        \register[21][8] ) );
  DFFRX1 \register_reg[21][7]  ( .D(n1740), .CK(clk), .RN(n2234), .Q(
        \register[21][7] ) );
  DFFRX1 \register_reg[21][6]  ( .D(n1741), .CK(clk), .RN(n2234), .Q(
        \register[21][6] ) );
  DFFRX1 \register_reg[21][5]  ( .D(n1742), .CK(clk), .RN(n2234), .Q(
        \register[21][5] ) );
  DFFRX1 \register_reg[21][4]  ( .D(n1743), .CK(clk), .RN(n2233), .Q(
        \register[21][4] ) );
  DFFRX1 \register_reg[25][8]  ( .D(n1867), .CK(clk), .RN(n2224), .Q(
        \register[25][8] ) );
  DFFRX1 \register_reg[25][7]  ( .D(n1868), .CK(clk), .RN(n2224), .Q(
        \register[25][7] ) );
  DFFRX1 \register_reg[25][6]  ( .D(n1869), .CK(clk), .RN(n2224), .Q(
        \register[25][6] ) );
  DFFRX1 \register_reg[25][5]  ( .D(n1870), .CK(clk), .RN(n2224), .Q(
        \register[25][5] ) );
  DFFRX1 \register_reg[25][4]  ( .D(n1871), .CK(clk), .RN(n2224), .Q(
        \register[25][4] ) );
  DFFRX1 \register_reg[29][8]  ( .D(n1995), .CK(clk), .RN(n2214), .Q(
        \register[29][8] ) );
  DFFRX1 \register_reg[29][7]  ( .D(n1996), .CK(clk), .RN(n2214), .Q(
        \register[29][7] ) );
  DFFRX1 \register_reg[29][6]  ( .D(n1997), .CK(clk), .RN(n2214), .Q(
        \register[29][6] ) );
  DFFRX1 \register_reg[29][5]  ( .D(n1998), .CK(clk), .RN(n2214), .Q(
        \register[29][5] ) );
  DFFRX1 \register_reg[29][4]  ( .D(n1999), .CK(clk), .RN(n2214), .Q(
        \register[29][4] ) );
  DFFRX1 \register_reg[1][3]  ( .D(n1104), .CK(clk), .RN(n2283), .Q(
        \register[1][3] ) );
  DFFRX1 \register_reg[1][2]  ( .D(n1105), .CK(clk), .RN(n2283), .Q(
        \register[1][2] ) );
  DFFRX1 \register_reg[1][1]  ( .D(n1106), .CK(clk), .RN(n2282), .Q(
        \register[1][1] ) );
  DFFRX1 \register_reg[1][0]  ( .D(n1107), .CK(clk), .RN(n2282), .Q(
        \register[1][0] ) );
  DFFRX1 \register_reg[5][3]  ( .D(n1232), .CK(clk), .RN(n2273), .Q(
        \register[5][3] ) );
  DFFRX1 \register_reg[5][2]  ( .D(n1233), .CK(clk), .RN(n2273), .Q(
        \register[5][2] ) );
  DFFRX1 \register_reg[5][1]  ( .D(n1234), .CK(clk), .RN(n2273), .Q(
        \register[5][1] ) );
  DFFRX1 \register_reg[5][0]  ( .D(n1235), .CK(clk), .RN(n2273), .Q(
        \register[5][0] ) );
  DFFRX1 \register_reg[9][3]  ( .D(n1360), .CK(clk), .RN(n2263), .Q(
        \register[9][3] ) );
  DFFRX1 \register_reg[9][2]  ( .D(n1361), .CK(clk), .RN(n2263), .Q(
        \register[9][2] ) );
  DFFRX1 \register_reg[9][1]  ( .D(n1362), .CK(clk), .RN(n2263), .Q(
        \register[9][1] ) );
  DFFRX1 \register_reg[9][0]  ( .D(n1363), .CK(clk), .RN(n2263), .Q(
        \register[9][0] ) );
  DFFRX1 \register_reg[13][3]  ( .D(n1488), .CK(clk), .RN(n2253), .Q(
        \register[13][3] ) );
  DFFRX1 \register_reg[13][2]  ( .D(n1489), .CK(clk), .RN(n2253), .Q(
        \register[13][2] ) );
  DFFRX1 \register_reg[13][1]  ( .D(n1490), .CK(clk), .RN(n2253), .Q(
        \register[13][1] ) );
  DFFRX1 \register_reg[13][0]  ( .D(n1491), .CK(clk), .RN(n2253), .Q(
        \register[13][0] ) );
  DFFRX1 \register_reg[17][3]  ( .D(n1616), .CK(clk), .RN(n2243), .Q(
        \register[17][3] ) );
  DFFRX1 \register_reg[17][2]  ( .D(n1617), .CK(clk), .RN(n2243), .Q(
        \register[17][2] ) );
  DFFRX1 \register_reg[17][1]  ( .D(n1618), .CK(clk), .RN(n2243), .Q(
        \register[17][1] ) );
  DFFRX1 \register_reg[17][0]  ( .D(n1619), .CK(clk), .RN(n2243), .Q(
        \register[17][0] ) );
  DFFRX1 \register_reg[21][3]  ( .D(n1744), .CK(clk), .RN(n2233), .Q(
        \register[21][3] ) );
  DFFRX1 \register_reg[21][2]  ( .D(n1745), .CK(clk), .RN(n2233), .Q(
        \register[21][2] ) );
  DFFRX1 \register_reg[21][1]  ( .D(n1746), .CK(clk), .RN(n2233), .Q(
        \register[21][1] ) );
  DFFRX1 \register_reg[21][0]  ( .D(n1747), .CK(clk), .RN(n2233), .Q(
        \register[21][0] ) );
  DFFRX1 \register_reg[25][3]  ( .D(n1872), .CK(clk), .RN(n2224), .Q(
        \register[25][3] ) );
  DFFRX1 \register_reg[25][2]  ( .D(n1873), .CK(clk), .RN(n2223), .Q(
        \register[25][2] ) );
  DFFRX1 \register_reg[25][0]  ( .D(n1875), .CK(clk), .RN(n2223), .Q(
        \register[25][0] ) );
  DFFRX1 \register_reg[29][3]  ( .D(n2000), .CK(clk), .RN(n2214), .Q(
        \register[29][3] ) );
  DFFRX1 \register_reg[29][1]  ( .D(n2002), .CK(clk), .RN(n2214), .Q(
        \register[29][1] ) );
  DFFRX1 \register_reg[29][2]  ( .D(n2001), .CK(clk), .RN(n2214), .Q(
        \register[29][2] ) );
  DFFRX1 \register_reg[0][8]  ( .D(n1067), .CK(clk), .RN(n2285), .Q(
        \register[0][8] ) );
  DFFRX1 \register_reg[0][7]  ( .D(n1068), .CK(clk), .RN(n2285), .Q(
        \register[0][7] ) );
  DFFRX1 \register_reg[0][6]  ( .D(n1069), .CK(clk), .RN(n2285), .Q(
        \register[0][6] ) );
  DFFRX1 \register_reg[0][5]  ( .D(n1070), .CK(clk), .RN(n2285), .Q(
        \register[0][5] ) );
  DFFRX1 \register_reg[0][4]  ( .D(n1071), .CK(clk), .RN(n2285), .Q(
        \register[0][4] ) );
  DFFRX1 \register_reg[4][8]  ( .D(n1195), .CK(clk), .RN(n2276), .Q(
        \register[4][8] ) );
  DFFRX1 \register_reg[4][7]  ( .D(n1196), .CK(clk), .RN(n2276), .Q(
        \register[4][7] ) );
  DFFRX1 \register_reg[4][6]  ( .D(n1197), .CK(clk), .RN(n2275), .Q(
        \register[4][6] ) );
  DFFRX1 \register_reg[4][5]  ( .D(n1198), .CK(clk), .RN(n2275), .Q(
        \register[4][5] ) );
  DFFRX1 \register_reg[4][4]  ( .D(n1199), .CK(clk), .RN(n2275), .Q(
        \register[4][4] ) );
  DFFRX1 \register_reg[8][8]  ( .D(n1323), .CK(clk), .RN(n2266), .Q(
        \register[8][8] ) );
  DFFRX1 \register_reg[8][7]  ( .D(n1324), .CK(clk), .RN(n2266), .Q(
        \register[8][7] ) );
  DFFRX1 \register_reg[8][6]  ( .D(n1325), .CK(clk), .RN(n2266), .Q(
        \register[8][6] ) );
  DFFRX1 \register_reg[8][5]  ( .D(n1326), .CK(clk), .RN(n2266), .Q(
        \register[8][5] ) );
  DFFRX1 \register_reg[8][4]  ( .D(n1327), .CK(clk), .RN(n2265), .Q(
        \register[8][4] ) );
  DFFRX1 \register_reg[12][8]  ( .D(n1451), .CK(clk), .RN(n2256), .Q(
        \register[12][8] ) );
  DFFRX1 \register_reg[12][7]  ( .D(n1452), .CK(clk), .RN(n2256), .Q(
        \register[12][7] ) );
  DFFRX1 \register_reg[12][6]  ( .D(n1453), .CK(clk), .RN(n2256), .Q(
        \register[12][6] ) );
  DFFRX1 \register_reg[12][5]  ( .D(n1454), .CK(clk), .RN(n2256), .Q(
        \register[12][5] ) );
  DFFRX1 \register_reg[12][4]  ( .D(n1455), .CK(clk), .RN(n2256), .Q(
        \register[12][4] ) );
  DFFRX1 \register_reg[16][8]  ( .D(n1579), .CK(clk), .RN(n2246), .Q(
        \register[16][8] ) );
  DFFRX1 \register_reg[16][7]  ( .D(n1580), .CK(clk), .RN(n2246), .Q(
        \register[16][7] ) );
  DFFRX1 \register_reg[16][6]  ( .D(n1581), .CK(clk), .RN(n2246), .Q(
        \register[16][6] ) );
  DFFRX1 \register_reg[16][5]  ( .D(n1582), .CK(clk), .RN(n2246), .Q(
        \register[16][5] ) );
  DFFRX1 \register_reg[16][4]  ( .D(n1583), .CK(clk), .RN(n2246), .Q(
        \register[16][4] ) );
  DFFRX1 \register_reg[20][8]  ( .D(n1707), .CK(clk), .RN(n2236), .Q(
        \register[20][8] ) );
  DFFRX1 \register_reg[20][7]  ( .D(n1708), .CK(clk), .RN(n2236), .Q(
        \register[20][7] ) );
  DFFRX1 \register_reg[20][6]  ( .D(n1709), .CK(clk), .RN(n2236), .Q(
        \register[20][6] ) );
  DFFRX1 \register_reg[20][5]  ( .D(n1710), .CK(clk), .RN(n2236), .Q(
        \register[20][5] ) );
  DFFRX1 \register_reg[20][4]  ( .D(n1711), .CK(clk), .RN(n2236), .Q(
        \register[20][4] ) );
  DFFRX1 \register_reg[24][8]  ( .D(n1835), .CK(clk), .RN(n2226), .Q(
        \register[24][8] ) );
  DFFRX1 \register_reg[24][7]  ( .D(n1836), .CK(clk), .RN(n2226), .Q(
        \register[24][7] ) );
  DFFRX1 \register_reg[24][6]  ( .D(n1837), .CK(clk), .RN(n2226), .Q(
        \register[24][6] ) );
  DFFRX1 \register_reg[24][5]  ( .D(n1838), .CK(clk), .RN(n2226), .Q(
        \register[24][5] ) );
  DFFRX1 \register_reg[24][4]  ( .D(n1839), .CK(clk), .RN(n2226), .Q(
        \register[24][4] ) );
  DFFRX1 \register_reg[28][8]  ( .D(n1963), .CK(clk), .RN(n2217), .Q(
        \register[28][8] ) );
  DFFRX1 \register_reg[28][7]  ( .D(n1964), .CK(clk), .RN(n2216), .Q(
        \register[28][7] ) );
  DFFRX1 \register_reg[28][6]  ( .D(n1965), .CK(clk), .RN(n2216), .Q(
        \register[28][6] ) );
  DFFRX1 \register_reg[28][5]  ( .D(n1966), .CK(clk), .RN(n2216), .Q(
        \register[28][5] ) );
  DFFRX1 \register_reg[28][4]  ( .D(n1967), .CK(clk), .RN(n2216), .Q(
        \register[28][4] ) );
  DFFRX1 \register_reg[0][3]  ( .D(n1072), .CK(clk), .RN(n2285), .Q(
        \register[0][3] ) );
  DFFRX1 \register_reg[0][2]  ( .D(n1073), .CK(clk), .RN(n2285), .Q(
        \register[0][2] ) );
  DFFRX1 \register_reg[0][1]  ( .D(n1074), .CK(clk), .RN(n2285), .Q(
        \register[0][1] ) );
  DFFRX1 \register_reg[0][0]  ( .D(n1075), .CK(clk), .RN(n2285), .Q(
        \register[0][0] ) );
  DFFRX1 \register_reg[4][3]  ( .D(n1200), .CK(clk), .RN(n2275), .Q(
        \register[4][3] ) );
  DFFRX1 \register_reg[4][2]  ( .D(n1201), .CK(clk), .RN(n2275), .Q(
        \register[4][2] ) );
  DFFRX1 \register_reg[4][1]  ( .D(n1202), .CK(clk), .RN(n2275), .Q(
        \register[4][1] ) );
  DFFRX1 \register_reg[4][0]  ( .D(n1203), .CK(clk), .RN(n2275), .Q(
        \register[4][0] ) );
  DFFRX1 \register_reg[8][3]  ( .D(n1328), .CK(clk), .RN(n2265), .Q(
        \register[8][3] ) );
  DFFRX1 \register_reg[8][2]  ( .D(n1329), .CK(clk), .RN(n2265), .Q(
        \register[8][2] ) );
  DFFRX1 \register_reg[8][1]  ( .D(n1330), .CK(clk), .RN(n2265), .Q(
        \register[8][1] ) );
  DFFRX1 \register_reg[8][0]  ( .D(n1331), .CK(clk), .RN(n2265), .Q(
        \register[8][0] ) );
  DFFRX1 \register_reg[12][3]  ( .D(n1456), .CK(clk), .RN(n2256), .Q(
        \register[12][3] ) );
  DFFRX1 \register_reg[12][2]  ( .D(n1457), .CK(clk), .RN(n2255), .Q(
        \register[12][2] ) );
  DFFRX1 \register_reg[12][1]  ( .D(n1458), .CK(clk), .RN(n2255), .Q(
        \register[12][1] ) );
  DFFRX1 \register_reg[12][0]  ( .D(n1459), .CK(clk), .RN(n2255), .Q(
        \register[12][0] ) );
  DFFRX1 \register_reg[16][3]  ( .D(n1584), .CK(clk), .RN(n2246), .Q(
        \register[16][3] ) );
  DFFRX1 \register_reg[16][2]  ( .D(n1585), .CK(clk), .RN(n2246), .Q(
        \register[16][2] ) );
  DFFRX1 \register_reg[16][1]  ( .D(n1586), .CK(clk), .RN(n2246), .Q(
        \register[16][1] ) );
  DFFRX1 \register_reg[16][0]  ( .D(n1587), .CK(clk), .RN(n2245), .Q(
        \register[16][0] ) );
  DFFRX1 \register_reg[20][3]  ( .D(n1712), .CK(clk), .RN(n2236), .Q(
        \register[20][3] ) );
  DFFRX1 \register_reg[20][2]  ( .D(n1713), .CK(clk), .RN(n2236), .Q(
        \register[20][2] ) );
  DFFRX1 \register_reg[20][1]  ( .D(n1714), .CK(clk), .RN(n2236), .Q(
        \register[20][1] ) );
  DFFRX1 \register_reg[24][3]  ( .D(n1840), .CK(clk), .RN(n2226), .Q(
        \register[24][3] ) );
  DFFRX1 \register_reg[24][2]  ( .D(n1841), .CK(clk), .RN(n2226), .Q(
        \register[24][2] ) );
  DFFRX1 \register_reg[24][1]  ( .D(n1842), .CK(clk), .RN(n2226), .Q(
        \register[24][1] ) );
  DFFRX1 \register_reg[24][0]  ( .D(n1843), .CK(clk), .RN(n2226), .Q(
        \register[24][0] ) );
  DFFRX1 \register_reg[28][3]  ( .D(n1968), .CK(clk), .RN(n2216), .Q(
        \register[28][3] ) );
  DFFRX1 \register_reg[28][1]  ( .D(n1970), .CK(clk), .RN(n2216), .Q(
        \register[28][1] ) );
  DFFRX1 \register_reg[28][2]  ( .D(n1969), .CK(clk), .RN(n2216), .Q(
        \register[28][2] ) );
  DFFRX1 \register_reg[2][8]  ( .D(n1131), .CK(clk), .RN(n2281), .Q(
        \register[2][8] ) );
  DFFRX1 \register_reg[2][7]  ( .D(n1132), .CK(clk), .RN(n2280), .Q(
        \register[2][7] ) );
  DFFRX1 \register_reg[2][6]  ( .D(n1133), .CK(clk), .RN(n2280), .Q(
        \register[2][6] ) );
  DFFRX1 \register_reg[2][5]  ( .D(n1134), .CK(clk), .RN(n2280), .Q(
        \register[2][5] ) );
  DFFRX1 \register_reg[2][4]  ( .D(n1135), .CK(clk), .RN(n2280), .Q(
        \register[2][4] ) );
  DFFRX1 \register_reg[6][8]  ( .D(n1259), .CK(clk), .RN(n2271), .Q(
        \register[6][8] ) );
  DFFRX1 \register_reg[6][7]  ( .D(n1260), .CK(clk), .RN(n2271), .Q(
        \register[6][7] ) );
  DFFRX1 \register_reg[6][6]  ( .D(n1261), .CK(clk), .RN(n2271), .Q(
        \register[6][6] ) );
  DFFRX1 \register_reg[6][5]  ( .D(n1262), .CK(clk), .RN(n2270), .Q(
        \register[6][5] ) );
  DFFRX1 \register_reg[6][4]  ( .D(n1263), .CK(clk), .RN(n2270), .Q(
        \register[6][4] ) );
  DFFRX1 \register_reg[10][8]  ( .D(n1387), .CK(clk), .RN(n2261), .Q(
        \register[10][8] ) );
  DFFRX1 \register_reg[10][7]  ( .D(n1388), .CK(clk), .RN(n2261), .Q(
        \register[10][7] ) );
  DFFRX1 \register_reg[10][6]  ( .D(n1389), .CK(clk), .RN(n2261), .Q(
        \register[10][6] ) );
  DFFRX1 \register_reg[10][5]  ( .D(n1390), .CK(clk), .RN(n2261), .Q(
        \register[10][5] ) );
  DFFRX1 \register_reg[10][4]  ( .D(n1391), .CK(clk), .RN(n2261), .Q(
        \register[10][4] ) );
  DFFRX1 \register_reg[14][8]  ( .D(n1515), .CK(clk), .RN(n2251), .Q(
        \register[14][8] ) );
  DFFRX1 \register_reg[14][7]  ( .D(n1516), .CK(clk), .RN(n2251), .Q(
        \register[14][7] ) );
  DFFRX1 \register_reg[14][6]  ( .D(n1517), .CK(clk), .RN(n2251), .Q(
        \register[14][6] ) );
  DFFRX1 \register_reg[14][5]  ( .D(n1518), .CK(clk), .RN(n2251), .Q(
        \register[14][5] ) );
  DFFRX1 \register_reg[14][4]  ( .D(n1519), .CK(clk), .RN(n2251), .Q(
        \register[14][4] ) );
  DFFRX1 \register_reg[18][8]  ( .D(n1643), .CK(clk), .RN(n2241), .Q(
        \register[18][8] ) );
  DFFRX1 \register_reg[18][7]  ( .D(n1644), .CK(clk), .RN(n2241), .Q(
        \register[18][7] ) );
  DFFRX1 \register_reg[18][6]  ( .D(n1645), .CK(clk), .RN(n2241), .Q(
        \register[18][6] ) );
  DFFRX1 \register_reg[18][5]  ( .D(n1646), .CK(clk), .RN(n2241), .Q(
        \register[18][5] ) );
  DFFRX1 \register_reg[18][4]  ( .D(n1647), .CK(clk), .RN(n2241), .Q(
        \register[18][4] ) );
  DFFRX1 \register_reg[22][8]  ( .D(n1771), .CK(clk), .RN(n2231), .Q(
        \register[22][8] ) );
  DFFRX1 \register_reg[22][7]  ( .D(n1772), .CK(clk), .RN(n2231), .Q(
        \register[22][7] ) );
  DFFRX1 \register_reg[22][6]  ( .D(n1773), .CK(clk), .RN(n2231), .Q(
        \register[22][6] ) );
  DFFRX1 \register_reg[22][5]  ( .D(n1774), .CK(clk), .RN(n2231), .Q(
        \register[22][5] ) );
  DFFRX1 \register_reg[22][4]  ( .D(n1775), .CK(clk), .RN(n2231), .Q(
        \register[22][4] ) );
  DFFRX1 \register_reg[26][8]  ( .D(n1899), .CK(clk), .RN(n2221), .Q(
        \register[26][8] ) );
  DFFRX1 \register_reg[26][7]  ( .D(n1900), .CK(clk), .RN(n2221), .Q(
        \register[26][7] ) );
  DFFRX1 \register_reg[26][6]  ( .D(n1901), .CK(clk), .RN(n2221), .Q(
        \register[26][6] ) );
  DFFRX1 \register_reg[26][5]  ( .D(n1902), .CK(clk), .RN(n2221), .Q(
        \register[26][5] ) );
  DFFRX1 \register_reg[26][4]  ( .D(n1903), .CK(clk), .RN(n2221), .Q(
        \register[26][4] ) );
  DFFRX1 \register_reg[30][8]  ( .D(n2027), .CK(clk), .RN(n2212), .Q(
        \register[30][8] ) );
  DFFRX1 \register_reg[30][7]  ( .D(n2028), .CK(clk), .RN(n2212), .Q(
        \register[30][7] ) );
  DFFRX1 \register_reg[30][6]  ( .D(n2029), .CK(clk), .RN(n2211), .Q(
        \register[30][6] ) );
  DFFRX1 \register_reg[30][5]  ( .D(n2030), .CK(clk), .RN(n2211), .Q(
        \register[30][5] ) );
  DFFRX1 \register_reg[30][4]  ( .D(n2031), .CK(clk), .RN(n2211), .Q(
        \register[30][4] ) );
  DFFRX1 \register_reg[2][3]  ( .D(n1136), .CK(clk), .RN(n2280), .Q(
        \register[2][3] ) );
  DFFRX1 \register_reg[2][2]  ( .D(n1137), .CK(clk), .RN(n2280), .Q(
        \register[2][2] ) );
  DFFRX1 \register_reg[2][1]  ( .D(n1138), .CK(clk), .RN(n2280), .Q(
        \register[2][1] ) );
  DFFRX1 \register_reg[2][0]  ( .D(n1139), .CK(clk), .RN(n2280), .Q(
        \register[2][0] ) );
  DFFRX1 \register_reg[6][3]  ( .D(n1264), .CK(clk), .RN(n2270), .Q(
        \register[6][3] ) );
  DFFRX1 \register_reg[6][2]  ( .D(n1265), .CK(clk), .RN(n2270), .Q(
        \register[6][2] ) );
  DFFRX1 \register_reg[6][1]  ( .D(n1266), .CK(clk), .RN(n2270), .Q(
        \register[6][1] ) );
  DFFRX1 \register_reg[6][0]  ( .D(n1267), .CK(clk), .RN(n2270), .Q(
        \register[6][0] ) );
  DFFRX1 \register_reg[10][3]  ( .D(n1392), .CK(clk), .RN(n2260), .Q(
        \register[10][3] ) );
  DFFRX1 \register_reg[10][2]  ( .D(n1393), .CK(clk), .RN(n2260), .Q(
        \register[10][2] ) );
  DFFRX1 \register_reg[10][1]  ( .D(n1394), .CK(clk), .RN(n2260), .Q(
        \register[10][1] ) );
  DFFRX1 \register_reg[10][0]  ( .D(n1395), .CK(clk), .RN(n2260), .Q(
        \register[10][0] ) );
  DFFRX1 \register_reg[14][3]  ( .D(n1520), .CK(clk), .RN(n2251), .Q(
        \register[14][3] ) );
  DFFRX1 \register_reg[14][2]  ( .D(n1521), .CK(clk), .RN(n2251), .Q(
        \register[14][2] ) );
  DFFRX1 \register_reg[14][1]  ( .D(n1522), .CK(clk), .RN(n2250), .Q(
        \register[14][1] ) );
  DFFRX1 \register_reg[14][0]  ( .D(n1523), .CK(clk), .RN(n2250), .Q(
        \register[14][0] ) );
  DFFRX1 \register_reg[18][3]  ( .D(n1648), .CK(clk), .RN(n2241), .Q(
        \register[18][3] ) );
  DFFRX1 \register_reg[18][2]  ( .D(n1649), .CK(clk), .RN(n2241), .Q(
        \register[18][2] ) );
  DFFRX1 \register_reg[18][1]  ( .D(n1650), .CK(clk), .RN(n2241), .Q(
        \register[18][1] ) );
  DFFRX1 \register_reg[18][0]  ( .D(n1651), .CK(clk), .RN(n2241), .Q(
        \register[18][0] ) );
  DFFRX1 \register_reg[22][3]  ( .D(n1776), .CK(clk), .RN(n2231), .Q(
        \register[22][3] ) );
  DFFRX1 \register_reg[22][2]  ( .D(n1777), .CK(clk), .RN(n2231), .Q(
        \register[22][2] ) );
  DFFRX1 \register_reg[22][1]  ( .D(n1778), .CK(clk), .RN(n2231), .Q(
        \register[22][1] ) );
  DFFRX1 \register_reg[22][0]  ( .D(n1779), .CK(clk), .RN(n2231), .Q(
        \register[22][0] ) );
  DFFRX1 \register_reg[26][3]  ( .D(n1904), .CK(clk), .RN(n2221), .Q(
        \register[26][3] ) );
  DFFRX1 \register_reg[26][2]  ( .D(n1905), .CK(clk), .RN(n2221), .Q(
        \register[26][2] ) );
  DFFRX1 \register_reg[26][1]  ( .D(n1906), .CK(clk), .RN(n2221), .Q(
        \register[26][1] ) );
  DFFRX1 \register_reg[26][0]  ( .D(n1907), .CK(clk), .RN(n2221), .Q(
        \register[26][0] ) );
  DFFRX1 \register_reg[30][3]  ( .D(n2032), .CK(clk), .RN(n2211), .Q(
        \register[30][3] ) );
  DFFRX1 \register_reg[30][1]  ( .D(n2034), .CK(clk), .RN(n2211), .Q(
        \register[30][1] ) );
  DFFRX1 \register_reg[30][2]  ( .D(n2033), .CK(clk), .RN(n2211), .Q(
        \register[30][2] ) );
  DFFRX1 \register_reg[25][1]  ( .D(n1874), .CK(clk), .RN(n2223), .Q(
        \register[25][1] ) );
  DFFRX1 \register_reg[29][0]  ( .D(n2003), .CK(clk), .RN(rst_n), .Q(
        \register[29][0] ), .QN(n2352) );
  DFFRX1 \register_reg[28][0]  ( .D(n1971), .CK(clk), .RN(n2216), .Q(
        \register[28][0] ), .QN(n2353) );
  DFFRX1 \register_reg[20][0]  ( .D(n1715), .CK(clk), .RN(n2236), .Q(
        \register[20][0] ) );
  DFFRX1 \register_reg[31][0]  ( .D(n2067), .CK(clk), .RN(n2209), .Q(
        \register[31][0] ), .QN(n65) );
  DFFRX1 \register_reg[30][0]  ( .D(n2035), .CK(clk), .RN(n2211), .Q(
        \register[30][0] ), .QN(n64) );
  MXI4X1 U3 ( .A(\register[28][0] ), .B(\register[29][0] ), .C(
        \register[30][0] ), .D(\register[31][0] ), .S0(n901), .S1(n858), .Y(
        n562) );
  MXI4X1 U4 ( .A(\register[16][0] ), .B(\register[17][0] ), .C(
        \register[18][0] ), .D(\register[19][0] ), .S0(n901), .S1(n858), .Y(
        n565) );
  MXI4X1 U5 ( .A(\register[24][0] ), .B(\register[25][0] ), .C(
        \register[26][0] ), .D(\register[27][0] ), .S0(n901), .S1(n858), .Y(
        n563) );
  MXI4X1 U6 ( .A(\register[0][0] ), .B(\register[1][0] ), .C(\register[2][0] ), 
        .D(\register[3][0] ), .S0(n902), .S1(n859), .Y(n569) );
  MXI4X1 U7 ( .A(\register[8][0] ), .B(\register[9][0] ), .C(\register[10][0] ), .D(\register[11][0] ), .S0(n902), .S1(n859), .Y(n567) );
  MXI4X1 U8 ( .A(\register[4][0] ), .B(\register[5][0] ), .C(\register[6][0] ), 
        .D(\register[7][0] ), .S0(n902), .S1(n859), .Y(n568) );
  MXI4X1 U9 ( .A(\register[20][1] ), .B(\register[21][1] ), .C(
        \register[22][1] ), .D(\register[23][1] ), .S0(n902), .S1(n859), .Y(
        n572) );
  MXI4X1 U10 ( .A(\register[16][1] ), .B(\register[17][1] ), .C(
        \register[18][1] ), .D(\register[19][1] ), .S0(n902), .S1(n859), .Y(
        n573) );
  MXI4X1 U11 ( .A(\register[28][1] ), .B(\register[29][1] ), .C(
        \register[30][1] ), .D(\register[31][1] ), .S0(n902), .S1(n859), .Y(
        n570) );
  MXI4X1 U12 ( .A(\register[0][1] ), .B(\register[1][1] ), .C(\register[2][1] ), .D(\register[3][1] ), .S0(n902), .S1(n859), .Y(n577) );
  MXI4X1 U13 ( .A(\register[8][1] ), .B(\register[9][1] ), .C(
        \register[10][1] ), .D(\register[11][1] ), .S0(n902), .S1(n859), .Y(
        n575) );
  MXI4X1 U14 ( .A(\register[4][1] ), .B(\register[5][1] ), .C(\register[6][1] ), .D(\register[7][1] ), .S0(n902), .S1(n859), .Y(n576) );
  MXI4X1 U15 ( .A(\register[0][14] ), .B(\register[1][14] ), .C(
        \register[2][14] ), .D(\register[3][14] ), .S0(n484), .S1(n443), .Y(
        n254) );
  MXI4X1 U16 ( .A(\register[0][16] ), .B(\register[1][16] ), .C(
        \register[2][16] ), .D(\register[3][16] ), .S0(n485), .S1(n444), .Y(
        n270) );
  MXI4X1 U17 ( .A(\register[0][17] ), .B(\register[1][17] ), .C(
        \register[2][17] ), .D(\register[3][17] ), .S0(n486), .S1(n445), .Y(
        n279) );
  MXI4X1 U18 ( .A(\register[0][24] ), .B(\register[1][24] ), .C(
        \register[2][24] ), .D(\register[3][24] ), .S0(n491), .S1(n450), .Y(
        n336) );
  MXI4X1 U19 ( .A(\register[0][25] ), .B(\register[1][25] ), .C(
        \register[2][25] ), .D(\register[3][25] ), .S0(n491), .S1(n450), .Y(
        n345) );
  CLKBUFX3 U20 ( .A(WriteData_i[31]), .Y(n2205) );
  MXI2X1 U21 ( .A(n82), .B(n83), .S0(n394), .Y(ReadData1_o[2]) );
  MXI2X1 U22 ( .A(n84), .B(n85), .S0(n394), .Y(ReadData1_o[3]) );
  MXI4X1 U23 ( .A(\register[0][22] ), .B(\register[1][22] ), .C(
        \register[2][22] ), .D(\register[3][22] ), .S0(n489), .S1(n448), .Y(
        n320) );
  MXI4X1 U24 ( .A(\register[0][1] ), .B(\register[1][1] ), .C(\register[2][1] ), .D(\register[3][1] ), .S0(n475), .S1(n434), .Y(n147) );
  MX4X1 U25 ( .A(n569), .B(n567), .C(n568), .D(n566), .S0(n824), .S1(n833), 
        .Y(n498) );
  MXI4X1 U26 ( .A(\register[12][0] ), .B(\register[13][0] ), .C(
        \register[14][0] ), .D(\register[15][0] ), .S0(n902), .S1(n859), .Y(
        n566) );
  MX4X1 U27 ( .A(n577), .B(n575), .C(n576), .D(n574), .S0(n824), .S1(n833), 
        .Y(n500) );
  MXI4X1 U28 ( .A(\register[12][1] ), .B(\register[13][1] ), .C(
        \register[14][1] ), .D(\register[15][1] ), .S0(n902), .S1(n859), .Y(
        n574) );
  MXI4X1 U29 ( .A(\register[24][3] ), .B(\register[25][3] ), .C(
        \register[26][3] ), .D(\register[27][3] ), .S0(n903), .S1(n860), .Y(
        n587) );
  NOR3X1 U30 ( .A(n2351), .B(n2350), .C(n1021), .Y(n1) );
  NOR3X1 U31 ( .A(n2351), .B(n2348), .C(n1021), .Y(n2) );
  NOR3X1 U32 ( .A(n2351), .B(n2347), .C(n1021), .Y(n3) );
  MXI4X1 U33 ( .A(\register[24][1] ), .B(\register[25][1] ), .C(
        \register[26][1] ), .D(\register[27][1] ), .S0(n902), .S1(n859), .Y(
        n571) );
  MXI4X1 U34 ( .A(\register[24][1] ), .B(\register[25][1] ), .C(
        \register[26][1] ), .D(\register[27][1] ), .S0(n475), .S1(n434), .Y(
        n141) );
  MXI2X1 U35 ( .A(n4), .B(n5), .S0(n394), .Y(ReadData1_o[1]) );
  BUFX2 U36 ( .A(n2203), .Y(n2201) );
  BUFX2 U37 ( .A(n2193), .Y(n2191) );
  BUFX2 U38 ( .A(n2198), .Y(n2196) );
  CLKBUFX3 U39 ( .A(n2178), .Y(n2176) );
  CLKBUFX3 U40 ( .A(n2183), .Y(n2181) );
  CLKBUFX3 U41 ( .A(n2188), .Y(n2186) );
  MXI4XL U42 ( .A(\register[0][0] ), .B(\register[1][0] ), .C(\register[2][0] ), .D(\register[3][0] ), .S0(n475), .S1(n434), .Y(n139) );
  MXI4XL U43 ( .A(\register[0][3] ), .B(\register[1][3] ), .C(\register[2][3] ), .D(\register[3][3] ), .S0(n477), .S1(n436), .Y(n163) );
  MXI4X1 U44 ( .A(\register[0][2] ), .B(\register[1][2] ), .C(\register[2][2] ), .D(\register[3][2] ), .S0(n476), .S1(n435), .Y(n155) );
  MXI4X1 U45 ( .A(\register[28][2] ), .B(\register[29][2] ), .C(
        \register[30][2] ), .D(\register[31][2] ), .S0(n903), .S1(n860), .Y(
        n578) );
  MXI4X1 U46 ( .A(\register[12][2] ), .B(\register[13][2] ), .C(
        \register[14][2] ), .D(\register[15][2] ), .S0(n903), .S1(n860), .Y(
        n582) );
  MXI4X1 U47 ( .A(\register[0][2] ), .B(\register[1][2] ), .C(\register[2][2] ), .D(\register[3][2] ), .S0(n903), .S1(n860), .Y(n585) );
  MXI4X1 U48 ( .A(\register[16][2] ), .B(\register[17][2] ), .C(
        \register[18][2] ), .D(\register[19][2] ), .S0(n903), .S1(n860), .Y(
        n581) );
  MXI4X1 U49 ( .A(\register[4][2] ), .B(\register[5][2] ), .C(\register[6][2] ), .D(\register[7][2] ), .S0(n903), .S1(n860), .Y(n584) );
  MXI4X1 U50 ( .A(\register[20][2] ), .B(\register[21][2] ), .C(
        \register[22][2] ), .D(\register[23][2] ), .S0(n903), .S1(n860), .Y(
        n580) );
  MXI4X1 U51 ( .A(\register[8][2] ), .B(\register[9][2] ), .C(
        \register[10][2] ), .D(\register[11][2] ), .S0(n903), .S1(n860), .Y(
        n583) );
  MXI4X1 U52 ( .A(\register[24][2] ), .B(\register[25][2] ), .C(
        \register[26][2] ), .D(\register[27][2] ), .S0(n903), .S1(n860), .Y(
        n579) );
  MXI4XL U53 ( .A(\register[16][0] ), .B(\register[17][0] ), .C(
        \register[18][0] ), .D(\register[19][0] ), .S0(n474), .S1(n433), .Y(
        n134) );
  MXI4XL U54 ( .A(\register[24][0] ), .B(\register[25][0] ), .C(
        \register[26][0] ), .D(\register[27][0] ), .S0(n474), .S1(n433), .Y(
        n132) );
  CLKBUFX2 U55 ( .A(n2203), .Y(n2202) );
  CLKBUFX2 U56 ( .A(n2198), .Y(n2197) );
  CLKBUFX2 U57 ( .A(n2193), .Y(n2192) );
  BUFX2 U58 ( .A(n2173), .Y(n2171) );
  BUFX2 U59 ( .A(n2168), .Y(n2166) );
  CLKBUFX2 U60 ( .A(n2188), .Y(n2187) );
  CLKBUFX2 U61 ( .A(n2183), .Y(n2182) );
  CLKBUFX2 U62 ( .A(n2178), .Y(n2177) );
  CLKBUFX2 U63 ( .A(n2173), .Y(n2172) );
  CLKBUFX2 U64 ( .A(n2168), .Y(n2167) );
  NOR2BX1 U65 ( .AN(n873), .B(Reg_W_i[2]), .Y(n70) );
  NOR2BX1 U66 ( .AN(n975), .B(Reg_W_i[2]), .Y(n172) );
  NOR2BX1 U67 ( .AN(n941), .B(Reg_W_i[2]), .Y(n138) );
  NOR2BX1 U68 ( .AN(n907), .B(Reg_W_i[2]), .Y(n104) );
  NOR2X1 U69 ( .A(Reg_W_i[3]), .B(Reg_W_i[4]), .Y(n69) );
  NOR2X1 U70 ( .A(n2355), .B(Reg_W_i[4]), .Y(n342) );
  MXI2X1 U71 ( .A(n96), .B(n97), .S0(n395), .Y(ReadData1_o[9]) );
  MXI2X1 U72 ( .A(n100), .B(n101), .S0(n395), .Y(ReadData1_o[11]) );
  MXI2X1 U73 ( .A(n92), .B(n93), .S0(n394), .Y(ReadData1_o[7]) );
  MXI2X1 U74 ( .A(n94), .B(n95), .S0(n395), .Y(ReadData1_o[8]) );
  MXI2X1 U75 ( .A(n98), .B(n99), .S0(n395), .Y(ReadData1_o[10]) );
  MXI2X1 U76 ( .A(n90), .B(n91), .S0(n394), .Y(ReadData1_o[6]) );
  MXI4XL U77 ( .A(\register[0][6] ), .B(\register[1][6] ), .C(\register[2][6] ), .D(\register[3][6] ), .S0(n479), .S1(n438), .Y(n188) );
  MXI2X1 U78 ( .A(n88), .B(n89), .S0(n394), .Y(ReadData1_o[5]) );
  MXI4XL U79 ( .A(\register[0][5] ), .B(\register[1][5] ), .C(\register[2][5] ), .D(\register[3][5] ), .S0(n478), .S1(n437), .Y(n180) );
  MXI2X1 U80 ( .A(n86), .B(n87), .S0(n394), .Y(ReadData1_o[4]) );
  MXI4XL U81 ( .A(\register[0][4] ), .B(\register[1][4] ), .C(\register[2][4] ), .D(\register[3][4] ), .S0(n477), .S1(n436), .Y(n171) );
  MXI2XL U82 ( .A(n504), .B(n505), .S0(n819), .Y(ReadData2_o[3]) );
  MXI4X2 U83 ( .A(\register[28][3] ), .B(\register[29][3] ), .C(
        \register[30][3] ), .D(\register[31][3] ), .S0(n903), .S1(n860), .Y(
        n586) );
  MXI2XL U84 ( .A(n506), .B(n507), .S0(n819), .Y(ReadData2_o[4]) );
  MXI2XL U85 ( .A(n508), .B(n509), .S0(n819), .Y(ReadData2_o[5]) );
  MXI2XL U86 ( .A(n510), .B(n511), .S0(n819), .Y(ReadData2_o[6]) );
  MX4X1 U87 ( .A(n147), .B(n145), .C(n146), .D(n144), .S0(n399), .S1(n408), 
        .Y(n4) );
  MX4X1 U88 ( .A(n143), .B(n141), .C(n142), .D(n140), .S0(n399), .S1(n408), 
        .Y(n5) );
  MXI4X2 U89 ( .A(\register[12][3] ), .B(\register[13][3] ), .C(
        \register[14][3] ), .D(\register[15][3] ), .S0(n904), .S1(n861), .Y(
        n590) );
  MXI4XL U90 ( .A(\register[28][3] ), .B(\register[29][3] ), .C(
        \register[30][3] ), .D(\register[31][3] ), .S0(n476), .S1(n435), .Y(
        n156) );
  MXI4XL U91 ( .A(\register[28][2] ), .B(\register[29][2] ), .C(
        \register[30][2] ), .D(\register[31][2] ), .S0(n476), .S1(n435), .Y(
        n148) );
  MXI4XL U92 ( .A(\register[12][3] ), .B(\register[13][3] ), .C(
        \register[14][3] ), .D(\register[15][3] ), .S0(n477), .S1(n436), .Y(
        n160) );
  MXI4XL U93 ( .A(\register[12][2] ), .B(\register[13][2] ), .C(
        \register[14][2] ), .D(\register[15][2] ), .S0(n476), .S1(n435), .Y(
        n152) );
  MXI4XL U94 ( .A(\register[28][5] ), .B(\register[29][5] ), .C(
        \register[30][5] ), .D(\register[31][5] ), .S0(n478), .S1(n437), .Y(
        n173) );
  MXI4XL U95 ( .A(\register[28][4] ), .B(\register[29][4] ), .C(
        \register[30][4] ), .D(\register[31][4] ), .S0(n477), .S1(n436), .Y(
        n164) );
  MXI4XL U96 ( .A(\register[12][5] ), .B(\register[13][5] ), .C(
        \register[14][5] ), .D(\register[15][5] ), .S0(n478), .S1(n437), .Y(
        n177) );
  MXI4XL U97 ( .A(\register[12][4] ), .B(\register[13][4] ), .C(
        \register[14][4] ), .D(\register[15][4] ), .S0(n477), .S1(n436), .Y(
        n168) );
  MXI4XL U98 ( .A(\register[28][6] ), .B(\register[29][6] ), .C(
        \register[30][6] ), .D(\register[31][6] ), .S0(n478), .S1(n437), .Y(
        n181) );
  MXI4XL U99 ( .A(\register[12][6] ), .B(\register[13][6] ), .C(
        \register[14][6] ), .D(\register[15][6] ), .S0(n479), .S1(n438), .Y(
        n185) );
  MXI4XL U100 ( .A(\register[12][0] ), .B(\register[13][0] ), .C(
        \register[14][0] ), .D(\register[15][0] ), .S0(n475), .S1(n434), .Y(
        n135) );
  MXI4X2 U101 ( .A(\register[0][3] ), .B(\register[1][3] ), .C(
        \register[2][3] ), .D(\register[3][3] ), .S0(n904), .S1(n861), .Y(n593) );
  MXI4X2 U102 ( .A(\register[16][3] ), .B(\register[17][3] ), .C(
        \register[18][3] ), .D(\register[19][3] ), .S0(n903), .S1(n860), .Y(
        n589) );
  MXI4XL U103 ( .A(\register[16][3] ), .B(\register[17][3] ), .C(
        \register[18][3] ), .D(\register[19][3] ), .S0(n476), .S1(n435), .Y(
        n159) );
  MXI4XL U104 ( .A(\register[16][2] ), .B(\register[17][2] ), .C(
        \register[18][2] ), .D(\register[19][2] ), .S0(n476), .S1(n435), .Y(
        n151) );
  MXI4XL U105 ( .A(\register[16][5] ), .B(\register[17][5] ), .C(
        \register[18][5] ), .D(\register[19][5] ), .S0(n478), .S1(n437), .Y(
        n176) );
  MXI4XL U106 ( .A(\register[16][4] ), .B(\register[17][4] ), .C(
        \register[18][4] ), .D(\register[19][4] ), .S0(n477), .S1(n436), .Y(
        n167) );
  MXI4XL U107 ( .A(\register[16][6] ), .B(\register[17][6] ), .C(
        \register[18][6] ), .D(\register[19][6] ), .S0(n478), .S1(n437), .Y(
        n184) );
  MXI4X2 U108 ( .A(\register[20][0] ), .B(\register[21][0] ), .C(
        \register[22][0] ), .D(\register[23][0] ), .S0(n901), .S1(n858), .Y(
        n564) );
  MXI4XL U109 ( .A(\register[20][0] ), .B(\register[21][0] ), .C(
        \register[22][0] ), .D(\register[23][0] ), .S0(n474), .S1(n433), .Y(
        n133) );
  MXI4X2 U110 ( .A(\register[4][3] ), .B(\register[5][3] ), .C(
        \register[6][3] ), .D(\register[7][3] ), .S0(n904), .S1(n861), .Y(n592) );
  MXI4X2 U111 ( .A(\register[20][3] ), .B(\register[21][3] ), .C(
        \register[22][3] ), .D(\register[23][3] ), .S0(n903), .S1(n860), .Y(
        n588) );
  MXI4XL U112 ( .A(\register[20][3] ), .B(\register[21][3] ), .C(
        \register[22][3] ), .D(\register[23][3] ), .S0(n476), .S1(n435), .Y(
        n158) );
  MXI4XL U113 ( .A(\register[20][2] ), .B(\register[21][2] ), .C(
        \register[22][2] ), .D(\register[23][2] ), .S0(n476), .S1(n435), .Y(
        n150) );
  MXI4XL U114 ( .A(\register[4][3] ), .B(\register[5][3] ), .C(
        \register[6][3] ), .D(\register[7][3] ), .S0(n477), .S1(n436), .Y(n162) );
  MXI4XL U115 ( .A(\register[4][2] ), .B(\register[5][2] ), .C(
        \register[6][2] ), .D(\register[7][2] ), .S0(n476), .S1(n435), .Y(n154) );
  MXI4XL U116 ( .A(\register[20][5] ), .B(\register[21][5] ), .C(
        \register[22][5] ), .D(\register[23][5] ), .S0(n478), .S1(n437), .Y(
        n175) );
  MXI4XL U117 ( .A(\register[20][4] ), .B(\register[21][4] ), .C(
        \register[22][4] ), .D(\register[23][4] ), .S0(n477), .S1(n436), .Y(
        n166) );
  MXI4XL U118 ( .A(\register[4][5] ), .B(\register[5][5] ), .C(
        \register[6][5] ), .D(\register[7][5] ), .S0(n478), .S1(n437), .Y(n179) );
  MXI4XL U119 ( .A(\register[4][4] ), .B(\register[5][4] ), .C(
        \register[6][4] ), .D(\register[7][4] ), .S0(n477), .S1(n436), .Y(n170) );
  MXI4XL U120 ( .A(\register[20][6] ), .B(\register[21][6] ), .C(
        \register[22][6] ), .D(\register[23][6] ), .S0(n478), .S1(n437), .Y(
        n183) );
  MXI4XL U121 ( .A(\register[4][6] ), .B(\register[5][6] ), .C(
        \register[6][6] ), .D(\register[7][6] ), .S0(n479), .S1(n438), .Y(n187) );
  MXI4XL U122 ( .A(\register[4][0] ), .B(\register[5][0] ), .C(
        \register[6][0] ), .D(\register[7][0] ), .S0(n475), .S1(n434), .Y(n137) );
  MXI4X2 U123 ( .A(\register[8][3] ), .B(\register[9][3] ), .C(
        \register[10][3] ), .D(\register[11][3] ), .S0(n904), .S1(n861), .Y(
        n591) );
  MXI4XL U124 ( .A(\register[24][3] ), .B(\register[25][3] ), .C(
        \register[26][3] ), .D(\register[27][3] ), .S0(n476), .S1(n435), .Y(
        n157) );
  MXI4XL U125 ( .A(\register[24][2] ), .B(\register[25][2] ), .C(
        \register[26][2] ), .D(\register[27][2] ), .S0(n476), .S1(n435), .Y(
        n149) );
  MXI4XL U126 ( .A(\register[8][3] ), .B(\register[9][3] ), .C(
        \register[10][3] ), .D(\register[11][3] ), .S0(n477), .S1(n436), .Y(
        n161) );
  MXI4XL U127 ( .A(\register[8][2] ), .B(\register[9][2] ), .C(
        \register[10][2] ), .D(\register[11][2] ), .S0(n476), .S1(n435), .Y(
        n153) );
  MXI4XL U128 ( .A(\register[24][5] ), .B(\register[25][5] ), .C(
        \register[26][5] ), .D(\register[27][5] ), .S0(n478), .S1(n437), .Y(
        n174) );
  MXI4XL U129 ( .A(\register[24][4] ), .B(\register[25][4] ), .C(
        \register[26][4] ), .D(\register[27][4] ), .S0(n477), .S1(n436), .Y(
        n165) );
  MXI4XL U130 ( .A(\register[8][5] ), .B(\register[9][5] ), .C(
        \register[10][5] ), .D(\register[11][5] ), .S0(n478), .S1(n437), .Y(
        n178) );
  MXI4XL U131 ( .A(\register[8][4] ), .B(\register[9][4] ), .C(
        \register[10][4] ), .D(\register[11][4] ), .S0(n477), .S1(n436), .Y(
        n169) );
  MXI4XL U132 ( .A(\register[24][6] ), .B(\register[25][6] ), .C(
        \register[26][6] ), .D(\register[27][6] ), .S0(n478), .S1(n437), .Y(
        n182) );
  MXI4XL U133 ( .A(\register[8][6] ), .B(\register[9][6] ), .C(
        \register[10][6] ), .D(\register[11][6] ), .S0(n479), .S1(n438), .Y(
        n186) );
  MXI4XL U134 ( .A(\register[8][0] ), .B(\register[9][0] ), .C(
        \register[10][0] ), .D(\register[11][0] ), .S0(n475), .S1(n434), .Y(
        n136) );
  MXI4XL U135 ( .A(\register[12][1] ), .B(\register[13][1] ), .C(
        \register[14][1] ), .D(\register[15][1] ), .S0(n475), .S1(n434), .Y(
        n144) );
  MXI4XL U136 ( .A(\register[28][1] ), .B(\register[29][1] ), .C(
        \register[30][1] ), .D(\register[31][1] ), .S0(n475), .S1(n434), .Y(
        n140) );
  MXI4XL U137 ( .A(\register[4][1] ), .B(\register[5][1] ), .C(
        \register[6][1] ), .D(\register[7][1] ), .S0(n475), .S1(n434), .Y(n146) );
  MXI4XL U138 ( .A(\register[20][1] ), .B(\register[21][1] ), .C(
        \register[22][1] ), .D(\register[23][1] ), .S0(n475), .S1(n434), .Y(
        n142) );
  MXI4XL U139 ( .A(\register[16][1] ), .B(\register[17][1] ), .C(
        \register[18][1] ), .D(\register[19][1] ), .S0(n475), .S1(n434), .Y(
        n143) );
  MXI4XL U140 ( .A(\register[8][1] ), .B(\register[9][1] ), .C(
        \register[10][1] ), .D(\register[11][1] ), .S0(n475), .S1(n434), .Y(
        n145) );
  MXI2X1 U141 ( .A(n105), .B(n106), .S0(n395), .Y(ReadData1_o[13]) );
  MXI2X1 U142 ( .A(n107), .B(n108), .S0(n395), .Y(ReadData1_o[15]) );
  MXI2X1 U143 ( .A(n102), .B(n103), .S0(n395), .Y(ReadData1_o[12]) );
  MXI2X1 U144 ( .A(n111), .B(n112), .S0(n395), .Y(ReadData1_o[19]) );
  MXI2X1 U145 ( .A(n109), .B(n110), .S0(n395), .Y(ReadData1_o[18]) );
  MX2XL U146 ( .A(\register[31][0] ), .B(n1026), .S0(n1025), .Y(n2067) );
  MX2XL U147 ( .A(\register[31][1] ), .B(n1031), .S0(n1025), .Y(n2066) );
  MX2XL U148 ( .A(\register[31][2] ), .B(n1036), .S0(n1025), .Y(n2065) );
  MX2XL U149 ( .A(\register[31][3] ), .B(n1041), .S0(n1025), .Y(n2064) );
  MX2XL U150 ( .A(\register[31][4] ), .B(n2070), .S0(n1025), .Y(n2063) );
  MX2XL U151 ( .A(\register[31][5] ), .B(n2075), .S0(n1025), .Y(n2062) );
  MX2XL U152 ( .A(\register[31][6] ), .B(n2080), .S0(n1025), .Y(n2061) );
  MX2XL U153 ( .A(\register[30][0] ), .B(n1026), .S0(n1020), .Y(n2035) );
  MX2XL U154 ( .A(\register[30][1] ), .B(n1031), .S0(n1020), .Y(n2034) );
  MX2XL U155 ( .A(\register[30][2] ), .B(n1036), .S0(n1020), .Y(n2033) );
  MX2XL U156 ( .A(\register[30][3] ), .B(n1041), .S0(n1020), .Y(n2032) );
  MX2XL U157 ( .A(\register[30][4] ), .B(n2070), .S0(n1020), .Y(n2031) );
  MX2XL U158 ( .A(\register[30][5] ), .B(n2075), .S0(n1020), .Y(n2030) );
  MX2XL U159 ( .A(\register[30][6] ), .B(n2080), .S0(n1020), .Y(n2029) );
  MX2XL U160 ( .A(\register[29][1] ), .B(n1031), .S0(n1017), .Y(n2002) );
  MX2XL U161 ( .A(\register[29][2] ), .B(n1036), .S0(n1017), .Y(n2001) );
  MX2XL U162 ( .A(\register[29][3] ), .B(n1041), .S0(n1017), .Y(n2000) );
  MX2XL U163 ( .A(\register[29][4] ), .B(n2070), .S0(n1017), .Y(n1999) );
  MX2XL U164 ( .A(\register[29][5] ), .B(n2075), .S0(n1017), .Y(n1998) );
  MX2XL U165 ( .A(\register[29][6] ), .B(n2080), .S0(n1017), .Y(n1997) );
  MX2XL U166 ( .A(\register[28][1] ), .B(n1031), .S0(n1014), .Y(n1970) );
  MX2XL U167 ( .A(\register[28][2] ), .B(n1036), .S0(n1014), .Y(n1969) );
  MX2XL U168 ( .A(\register[28][3] ), .B(n1041), .S0(n1014), .Y(n1968) );
  MX2XL U169 ( .A(\register[28][4] ), .B(n2070), .S0(n1014), .Y(n1967) );
  MX2XL U170 ( .A(\register[28][5] ), .B(n2075), .S0(n1014), .Y(n1966) );
  MX2XL U171 ( .A(\register[28][6] ), .B(n2080), .S0(n1014), .Y(n1965) );
  MX2XL U172 ( .A(\register[27][0] ), .B(n1026), .S0(n1011), .Y(n1939) );
  MX2XL U173 ( .A(\register[27][1] ), .B(n1031), .S0(n1011), .Y(n1938) );
  MX2XL U174 ( .A(\register[27][2] ), .B(n1036), .S0(n1011), .Y(n1937) );
  MX2XL U175 ( .A(\register[27][3] ), .B(n1041), .S0(n1011), .Y(n1936) );
  MX2XL U176 ( .A(\register[27][4] ), .B(n2070), .S0(n1011), .Y(n1935) );
  MX2XL U177 ( .A(\register[27][5] ), .B(n2075), .S0(n1011), .Y(n1934) );
  MX2XL U178 ( .A(\register[27][6] ), .B(n2080), .S0(n1011), .Y(n1933) );
  MX2XL U179 ( .A(\register[26][0] ), .B(n1026), .S0(n1008), .Y(n1907) );
  MX2XL U180 ( .A(\register[26][1] ), .B(n1031), .S0(n1008), .Y(n1906) );
  MX2XL U181 ( .A(\register[26][2] ), .B(n1036), .S0(n1008), .Y(n1905) );
  MX2XL U182 ( .A(\register[26][3] ), .B(n1041), .S0(n1008), .Y(n1904) );
  MX2XL U183 ( .A(\register[26][4] ), .B(n2070), .S0(n1008), .Y(n1903) );
  MX2XL U184 ( .A(\register[26][5] ), .B(n2075), .S0(n1008), .Y(n1902) );
  MX2XL U185 ( .A(\register[26][6] ), .B(n2080), .S0(n1008), .Y(n1901) );
  MX2XL U186 ( .A(\register[25][0] ), .B(n1026), .S0(n1005), .Y(n1875) );
  MX2XL U187 ( .A(\register[25][1] ), .B(n1031), .S0(n1005), .Y(n1874) );
  MX2XL U188 ( .A(\register[25][2] ), .B(n1036), .S0(n1005), .Y(n1873) );
  MX2XL U189 ( .A(\register[25][3] ), .B(n1041), .S0(n1005), .Y(n1872) );
  MX2XL U190 ( .A(\register[25][4] ), .B(n2070), .S0(n1005), .Y(n1871) );
  MX2XL U191 ( .A(\register[25][5] ), .B(n2075), .S0(n1005), .Y(n1870) );
  MX2XL U192 ( .A(\register[25][6] ), .B(n2080), .S0(n1005), .Y(n1869) );
  MX2XL U193 ( .A(\register[24][0] ), .B(n1026), .S0(n1002), .Y(n1843) );
  MX2XL U194 ( .A(\register[24][1] ), .B(n1031), .S0(n1002), .Y(n1842) );
  MX2XL U195 ( .A(\register[24][2] ), .B(n1036), .S0(n1002), .Y(n1841) );
  MX2XL U196 ( .A(\register[24][3] ), .B(n1041), .S0(n1002), .Y(n1840) );
  MX2XL U197 ( .A(\register[24][4] ), .B(n2070), .S0(n1002), .Y(n1839) );
  MX2XL U198 ( .A(\register[24][5] ), .B(n2075), .S0(n1002), .Y(n1838) );
  MX2XL U199 ( .A(\register[24][6] ), .B(n2080), .S0(n1002), .Y(n1837) );
  MX2XL U200 ( .A(\register[23][0] ), .B(n1026), .S0(n999), .Y(n1811) );
  MX2XL U201 ( .A(\register[23][1] ), .B(n1031), .S0(n999), .Y(n1810) );
  MX2XL U202 ( .A(\register[23][2] ), .B(n1036), .S0(n999), .Y(n1809) );
  MX2XL U203 ( .A(\register[23][3] ), .B(n1041), .S0(n999), .Y(n1808) );
  MX2XL U204 ( .A(\register[23][4] ), .B(n2070), .S0(n999), .Y(n1807) );
  MX2XL U205 ( .A(\register[23][5] ), .B(n2075), .S0(n999), .Y(n1806) );
  MX2XL U206 ( .A(\register[23][6] ), .B(n2080), .S0(n999), .Y(n1805) );
  MX2XL U207 ( .A(\register[22][0] ), .B(n1026), .S0(n996), .Y(n1779) );
  MX2XL U208 ( .A(\register[22][1] ), .B(n1031), .S0(n996), .Y(n1778) );
  MX2XL U209 ( .A(\register[22][2] ), .B(n1036), .S0(n996), .Y(n1777) );
  MX2XL U210 ( .A(\register[22][3] ), .B(n1041), .S0(n996), .Y(n1776) );
  MX2XL U211 ( .A(\register[22][4] ), .B(n2070), .S0(n996), .Y(n1775) );
  MX2XL U212 ( .A(\register[22][5] ), .B(n2075), .S0(n996), .Y(n1774) );
  MX2XL U213 ( .A(\register[22][6] ), .B(n2080), .S0(n996), .Y(n1773) );
  MX2XL U214 ( .A(\register[21][0] ), .B(n1026), .S0(n993), .Y(n1747) );
  MX2XL U215 ( .A(\register[21][1] ), .B(n1031), .S0(n993), .Y(n1746) );
  MX2XL U216 ( .A(\register[21][2] ), .B(n1036), .S0(n993), .Y(n1745) );
  MX2XL U217 ( .A(\register[21][3] ), .B(n1041), .S0(n993), .Y(n1744) );
  MX2XL U218 ( .A(\register[21][4] ), .B(n2070), .S0(n993), .Y(n1743) );
  MX2XL U219 ( .A(\register[21][5] ), .B(n2075), .S0(n993), .Y(n1742) );
  MX2XL U220 ( .A(\register[21][6] ), .B(n2080), .S0(n993), .Y(n1741) );
  MX2XL U221 ( .A(\register[20][1] ), .B(n1031), .S0(n990), .Y(n1714) );
  MX2XL U222 ( .A(\register[20][2] ), .B(n1036), .S0(n990), .Y(n1713) );
  MX2XL U223 ( .A(\register[20][3] ), .B(n1041), .S0(n990), .Y(n1712) );
  MX2XL U224 ( .A(\register[20][4] ), .B(n2070), .S0(n990), .Y(n1711) );
  MX2XL U225 ( .A(\register[20][5] ), .B(n2075), .S0(n990), .Y(n1710) );
  MX2XL U226 ( .A(\register[20][6] ), .B(n2080), .S0(n990), .Y(n1709) );
  MX2XL U227 ( .A(\register[19][0] ), .B(n1027), .S0(n987), .Y(n1683) );
  MX2XL U228 ( .A(\register[19][1] ), .B(n1032), .S0(n987), .Y(n1682) );
  MX2XL U229 ( .A(\register[19][2] ), .B(n1037), .S0(n987), .Y(n1681) );
  MX2XL U230 ( .A(\register[19][3] ), .B(n1042), .S0(n987), .Y(n1680) );
  MX2XL U231 ( .A(\register[19][4] ), .B(n2071), .S0(n987), .Y(n1679) );
  MX2XL U232 ( .A(\register[19][5] ), .B(n2076), .S0(n987), .Y(n1678) );
  MX2XL U233 ( .A(\register[19][6] ), .B(n2081), .S0(n987), .Y(n1677) );
  MX2XL U234 ( .A(\register[18][0] ), .B(n1027), .S0(n984), .Y(n1651) );
  MX2XL U235 ( .A(\register[18][1] ), .B(n1032), .S0(n984), .Y(n1650) );
  MX2XL U236 ( .A(\register[18][2] ), .B(n1037), .S0(n984), .Y(n1649) );
  MX2XL U237 ( .A(\register[18][3] ), .B(n1042), .S0(n984), .Y(n1648) );
  MX2XL U238 ( .A(\register[18][4] ), .B(n2071), .S0(n984), .Y(n1647) );
  MX2XL U239 ( .A(\register[18][5] ), .B(n2076), .S0(n984), .Y(n1646) );
  MX2XL U240 ( .A(\register[18][6] ), .B(n2081), .S0(n984), .Y(n1645) );
  MX2XL U241 ( .A(\register[17][0] ), .B(n1027), .S0(n981), .Y(n1619) );
  MX2XL U242 ( .A(\register[17][1] ), .B(n1032), .S0(n981), .Y(n1618) );
  MX2XL U243 ( .A(\register[17][2] ), .B(n1037), .S0(n981), .Y(n1617) );
  MX2XL U244 ( .A(\register[17][3] ), .B(n1042), .S0(n981), .Y(n1616) );
  MX2XL U245 ( .A(\register[17][4] ), .B(n2071), .S0(n981), .Y(n1615) );
  MX2XL U246 ( .A(\register[17][5] ), .B(n2076), .S0(n981), .Y(n1614) );
  MX2XL U247 ( .A(\register[17][6] ), .B(n2081), .S0(n981), .Y(n1613) );
  MX2XL U248 ( .A(\register[16][0] ), .B(n1027), .S0(n978), .Y(n1587) );
  MX2XL U249 ( .A(\register[16][1] ), .B(n1032), .S0(n978), .Y(n1586) );
  MX2XL U250 ( .A(\register[16][2] ), .B(n1037), .S0(n978), .Y(n1585) );
  MX2XL U251 ( .A(\register[16][3] ), .B(n1042), .S0(n978), .Y(n1584) );
  MX2XL U252 ( .A(\register[16][4] ), .B(n2071), .S0(n978), .Y(n1583) );
  MX2XL U253 ( .A(\register[16][5] ), .B(n2076), .S0(n978), .Y(n1582) );
  MX2XL U254 ( .A(\register[16][6] ), .B(n2081), .S0(n978), .Y(n1581) );
  MX2XL U255 ( .A(\register[15][0] ), .B(n1027), .S0(n974), .Y(n1555) );
  MX2XL U256 ( .A(\register[15][1] ), .B(n1032), .S0(n974), .Y(n1554) );
  MX2XL U257 ( .A(\register[15][2] ), .B(n1037), .S0(n974), .Y(n1553) );
  MX2XL U258 ( .A(\register[15][3] ), .B(n1042), .S0(n974), .Y(n1552) );
  MX2XL U259 ( .A(\register[15][4] ), .B(n2071), .S0(n974), .Y(n1551) );
  MX2XL U260 ( .A(\register[15][5] ), .B(n2076), .S0(n974), .Y(n1550) );
  MX2XL U261 ( .A(\register[15][6] ), .B(n2081), .S0(n974), .Y(n1549) );
  MX2XL U262 ( .A(\register[14][0] ), .B(n1027), .S0(n971), .Y(n1523) );
  MX2XL U263 ( .A(\register[14][1] ), .B(n1032), .S0(n971), .Y(n1522) );
  MX2XL U264 ( .A(\register[14][2] ), .B(n1037), .S0(n971), .Y(n1521) );
  MX2XL U265 ( .A(\register[14][3] ), .B(n1042), .S0(n971), .Y(n1520) );
  MX2XL U266 ( .A(\register[14][4] ), .B(n2071), .S0(n971), .Y(n1519) );
  MX2XL U267 ( .A(\register[14][5] ), .B(n2076), .S0(n971), .Y(n1518) );
  MX2XL U268 ( .A(\register[14][6] ), .B(n2081), .S0(n971), .Y(n1517) );
  MX2XL U269 ( .A(\register[13][0] ), .B(n1027), .S0(n968), .Y(n1491) );
  MX2XL U270 ( .A(\register[13][1] ), .B(n1032), .S0(n968), .Y(n1490) );
  MX2XL U271 ( .A(\register[13][2] ), .B(n1037), .S0(n968), .Y(n1489) );
  MX2XL U272 ( .A(\register[13][3] ), .B(n1042), .S0(n968), .Y(n1488) );
  MX2XL U273 ( .A(\register[13][4] ), .B(n2071), .S0(n968), .Y(n1487) );
  MX2XL U274 ( .A(\register[13][5] ), .B(n2076), .S0(n968), .Y(n1486) );
  MX2XL U275 ( .A(\register[13][6] ), .B(n2081), .S0(n968), .Y(n1485) );
  MX2XL U276 ( .A(\register[12][0] ), .B(n1027), .S0(n965), .Y(n1459) );
  MX2XL U277 ( .A(\register[12][1] ), .B(n1032), .S0(n965), .Y(n1458) );
  MX2XL U278 ( .A(\register[12][2] ), .B(n1037), .S0(n965), .Y(n1457) );
  MX2XL U279 ( .A(\register[12][3] ), .B(n1042), .S0(n965), .Y(n1456) );
  MX2XL U280 ( .A(\register[12][4] ), .B(n2071), .S0(n965), .Y(n1455) );
  MX2XL U281 ( .A(\register[12][5] ), .B(n2076), .S0(n965), .Y(n1454) );
  MX2XL U282 ( .A(\register[12][6] ), .B(n2081), .S0(n965), .Y(n1453) );
  MX2XL U283 ( .A(\register[11][0] ), .B(n1027), .S0(n962), .Y(n1427) );
  MX2XL U284 ( .A(\register[11][1] ), .B(n1032), .S0(n962), .Y(n1426) );
  MX2XL U285 ( .A(\register[11][2] ), .B(n1037), .S0(n962), .Y(n1425) );
  MX2XL U286 ( .A(\register[11][3] ), .B(n1042), .S0(n962), .Y(n1424) );
  MX2XL U287 ( .A(\register[11][4] ), .B(n2071), .S0(n962), .Y(n1423) );
  MX2XL U288 ( .A(\register[11][5] ), .B(n2076), .S0(n962), .Y(n1422) );
  MX2XL U289 ( .A(\register[11][6] ), .B(n2081), .S0(n962), .Y(n1421) );
  MX2XL U290 ( .A(\register[10][0] ), .B(n1027), .S0(n959), .Y(n1395) );
  MX2XL U291 ( .A(\register[10][1] ), .B(n1032), .S0(n959), .Y(n1394) );
  MX2XL U292 ( .A(\register[10][2] ), .B(n1037), .S0(n959), .Y(n1393) );
  MX2XL U293 ( .A(\register[10][3] ), .B(n1042), .S0(n959), .Y(n1392) );
  MX2XL U294 ( .A(\register[10][4] ), .B(n2071), .S0(n959), .Y(n1391) );
  MX2XL U295 ( .A(\register[10][5] ), .B(n2076), .S0(n959), .Y(n1390) );
  MX2XL U296 ( .A(\register[10][6] ), .B(n2081), .S0(n959), .Y(n1389) );
  MX2XL U297 ( .A(\register[9][0] ), .B(n1027), .S0(n956), .Y(n1363) );
  MX2XL U298 ( .A(\register[9][1] ), .B(n1032), .S0(n956), .Y(n1362) );
  MX2XL U299 ( .A(\register[9][2] ), .B(n1037), .S0(n956), .Y(n1361) );
  MX2XL U300 ( .A(\register[9][3] ), .B(n1042), .S0(n956), .Y(n1360) );
  MX2XL U301 ( .A(\register[9][4] ), .B(n2071), .S0(n956), .Y(n1359) );
  MX2XL U302 ( .A(\register[9][5] ), .B(n2076), .S0(n956), .Y(n1358) );
  MX2XL U303 ( .A(\register[9][6] ), .B(n2081), .S0(n956), .Y(n1357) );
  MX2XL U304 ( .A(\register[8][0] ), .B(n1027), .S0(n953), .Y(n1331) );
  MX2XL U305 ( .A(\register[8][1] ), .B(n1032), .S0(n953), .Y(n1330) );
  MX2XL U306 ( .A(\register[8][2] ), .B(n1037), .S0(n953), .Y(n1329) );
  MX2XL U307 ( .A(\register[8][3] ), .B(n1042), .S0(n953), .Y(n1328) );
  MX2XL U308 ( .A(\register[8][4] ), .B(n2071), .S0(n953), .Y(n1327) );
  MX2XL U309 ( .A(\register[8][5] ), .B(n2076), .S0(n953), .Y(n1326) );
  MX2XL U310 ( .A(\register[8][6] ), .B(n2081), .S0(n953), .Y(n1325) );
  MX2XL U311 ( .A(\register[7][0] ), .B(n1028), .S0(n950), .Y(n1299) );
  MX2XL U312 ( .A(\register[7][1] ), .B(n1033), .S0(n950), .Y(n1298) );
  MX2XL U313 ( .A(\register[7][2] ), .B(n1038), .S0(n950), .Y(n1297) );
  MX2XL U314 ( .A(\register[7][3] ), .B(n1043), .S0(n950), .Y(n1296) );
  MX2XL U315 ( .A(\register[7][4] ), .B(n2072), .S0(n950), .Y(n1295) );
  MX2XL U316 ( .A(\register[7][5] ), .B(n2077), .S0(n950), .Y(n1294) );
  MX2XL U317 ( .A(\register[7][6] ), .B(n2082), .S0(n950), .Y(n1293) );
  MX2XL U318 ( .A(\register[6][0] ), .B(n1028), .S0(n947), .Y(n1267) );
  MX2XL U319 ( .A(\register[6][1] ), .B(n1033), .S0(n947), .Y(n1266) );
  MX2XL U320 ( .A(\register[6][2] ), .B(n1038), .S0(n947), .Y(n1265) );
  MX2XL U321 ( .A(\register[6][3] ), .B(n1043), .S0(n947), .Y(n1264) );
  MX2XL U322 ( .A(\register[6][4] ), .B(n2072), .S0(n947), .Y(n1263) );
  MX2XL U323 ( .A(\register[6][5] ), .B(n2077), .S0(n947), .Y(n1262) );
  MX2XL U324 ( .A(\register[6][6] ), .B(n2082), .S0(n947), .Y(n1261) );
  MX2XL U325 ( .A(\register[5][0] ), .B(n1028), .S0(n944), .Y(n1235) );
  MX2XL U326 ( .A(\register[5][1] ), .B(n1033), .S0(n944), .Y(n1234) );
  MX2XL U327 ( .A(\register[5][2] ), .B(n1038), .S0(n944), .Y(n1233) );
  MX2XL U328 ( .A(\register[5][3] ), .B(n1043), .S0(n944), .Y(n1232) );
  MX2XL U329 ( .A(\register[5][4] ), .B(n2072), .S0(n944), .Y(n1231) );
  MX2XL U330 ( .A(\register[5][5] ), .B(n2077), .S0(n944), .Y(n1230) );
  MX2XL U331 ( .A(\register[5][6] ), .B(n2082), .S0(n944), .Y(n1229) );
  MX2XL U332 ( .A(\register[4][0] ), .B(n1028), .S0(n940), .Y(n1203) );
  MX2XL U333 ( .A(\register[4][1] ), .B(n1033), .S0(n940), .Y(n1202) );
  MX2XL U334 ( .A(\register[4][2] ), .B(n1038), .S0(n940), .Y(n1201) );
  MX2XL U335 ( .A(\register[4][3] ), .B(n1043), .S0(n940), .Y(n1200) );
  MX2XL U336 ( .A(\register[4][4] ), .B(n2072), .S0(n940), .Y(n1199) );
  MX2XL U337 ( .A(\register[4][5] ), .B(n2077), .S0(n940), .Y(n1198) );
  MX2XL U338 ( .A(\register[4][6] ), .B(n2082), .S0(n940), .Y(n1197) );
  MX2XL U339 ( .A(\register[3][0] ), .B(n1028), .S0(n937), .Y(n1171) );
  MX2XL U340 ( .A(\register[3][1] ), .B(n1033), .S0(n937), .Y(n1170) );
  MX2XL U341 ( .A(\register[3][2] ), .B(n1038), .S0(n937), .Y(n1169) );
  MX2XL U342 ( .A(\register[3][3] ), .B(n1043), .S0(n937), .Y(n1168) );
  MX2XL U343 ( .A(\register[3][4] ), .B(n2072), .S0(n937), .Y(n1167) );
  MX2XL U344 ( .A(\register[3][5] ), .B(n2077), .S0(n937), .Y(n1166) );
  MX2XL U345 ( .A(\register[3][6] ), .B(n2082), .S0(n937), .Y(n1165) );
  MX2XL U346 ( .A(\register[2][0] ), .B(n1028), .S0(n934), .Y(n1139) );
  MX2XL U347 ( .A(\register[2][1] ), .B(n1033), .S0(n934), .Y(n1138) );
  MX2XL U348 ( .A(\register[2][2] ), .B(n1038), .S0(n934), .Y(n1137) );
  MX2XL U349 ( .A(\register[2][3] ), .B(n1043), .S0(n934), .Y(n1136) );
  MX2XL U350 ( .A(\register[2][4] ), .B(n2072), .S0(n934), .Y(n1135) );
  MX2XL U351 ( .A(\register[2][5] ), .B(n2077), .S0(n934), .Y(n1134) );
  MX2XL U352 ( .A(\register[2][6] ), .B(n2082), .S0(n934), .Y(n1133) );
  MX2XL U353 ( .A(\register[1][0] ), .B(n1028), .S0(n931), .Y(n1107) );
  MX2XL U354 ( .A(\register[1][1] ), .B(n1033), .S0(n931), .Y(n1106) );
  MX2XL U355 ( .A(\register[1][2] ), .B(n1038), .S0(n931), .Y(n1105) );
  MX2XL U356 ( .A(\register[1][3] ), .B(n1043), .S0(n931), .Y(n1104) );
  MX2XL U357 ( .A(\register[1][4] ), .B(n2072), .S0(n931), .Y(n1103) );
  MX2XL U358 ( .A(\register[1][5] ), .B(n2077), .S0(n931), .Y(n1102) );
  MX2XL U359 ( .A(\register[1][6] ), .B(n2082), .S0(n931), .Y(n1101) );
  MX2XL U360 ( .A(\register[0][0] ), .B(n1028), .S0(n928), .Y(n1075) );
  MX2XL U361 ( .A(\register[0][1] ), .B(n1033), .S0(n928), .Y(n1074) );
  MX2XL U362 ( .A(\register[0][2] ), .B(n1038), .S0(n928), .Y(n1073) );
  MX2XL U363 ( .A(\register[0][3] ), .B(n1043), .S0(n928), .Y(n1072) );
  MX2XL U364 ( .A(\register[0][4] ), .B(n2072), .S0(n928), .Y(n1071) );
  MX2XL U365 ( .A(\register[0][5] ), .B(n2077), .S0(n928), .Y(n1070) );
  MX2XL U366 ( .A(\register[0][6] ), .B(n2082), .S0(n928), .Y(n1069) );
  MXI2X1 U367 ( .A(n115), .B(n116), .S0(n396), .Y(ReadData1_o[21]) );
  MXI2X1 U368 ( .A(n119), .B(n120), .S0(n396), .Y(ReadData1_o[26]) );
  MXI2X1 U369 ( .A(n113), .B(n114), .S0(n396), .Y(ReadData1_o[20]) );
  MXI2X1 U370 ( .A(n117), .B(n118), .S0(n396), .Y(ReadData1_o[23]) );
  MXI2X1 U371 ( .A(n121), .B(n122), .S0(n396), .Y(ReadData1_o[27]) );
  MXI2X1 U372 ( .A(n125), .B(n126), .S0(n396), .Y(ReadData1_o[29]) );
  MXI2X1 U373 ( .A(n123), .B(n124), .S0(n396), .Y(ReadData1_o[28]) );
  CLKBUFX3 U374 ( .A(n2321), .Y(n2220) );
  CLKBUFX3 U375 ( .A(n2321), .Y(n2221) );
  CLKBUFX3 U376 ( .A(n2320), .Y(n2222) );
  CLKBUFX3 U377 ( .A(n2320), .Y(n2223) );
  CLKBUFX3 U378 ( .A(n2319), .Y(n2224) );
  CLKBUFX3 U379 ( .A(n2319), .Y(n2225) );
  CLKBUFX3 U380 ( .A(n2318), .Y(n2226) );
  CLKBUFX3 U381 ( .A(n2318), .Y(n2227) );
  CLKBUFX3 U382 ( .A(n2317), .Y(n2228) );
  CLKBUFX3 U383 ( .A(n2317), .Y(n2229) );
  CLKBUFX3 U384 ( .A(n2316), .Y(n2230) );
  CLKBUFX3 U385 ( .A(n2316), .Y(n2231) );
  CLKBUFX3 U386 ( .A(n2315), .Y(n2232) );
  CLKBUFX3 U387 ( .A(n2315), .Y(n2233) );
  CLKBUFX3 U388 ( .A(n2314), .Y(n2234) );
  CLKBUFX3 U389 ( .A(n2314), .Y(n2235) );
  CLKBUFX3 U390 ( .A(n2313), .Y(n2236) );
  CLKBUFX3 U391 ( .A(n2313), .Y(n2237) );
  CLKBUFX3 U392 ( .A(n2312), .Y(n2238) );
  CLKBUFX3 U393 ( .A(n2312), .Y(n2239) );
  CLKBUFX3 U394 ( .A(n2311), .Y(n2240) );
  CLKBUFX3 U395 ( .A(n2311), .Y(n2241) );
  CLKBUFX3 U396 ( .A(n2310), .Y(n2242) );
  CLKBUFX3 U397 ( .A(n2310), .Y(n2243) );
  CLKBUFX3 U398 ( .A(n2309), .Y(n2244) );
  CLKBUFX3 U399 ( .A(n2309), .Y(n2245) );
  CLKBUFX3 U400 ( .A(n2308), .Y(n2246) );
  CLKBUFX3 U401 ( .A(n2308), .Y(n2247) );
  CLKBUFX3 U402 ( .A(n2307), .Y(n2248) );
  CLKBUFX3 U403 ( .A(n2307), .Y(n2249) );
  CLKBUFX3 U404 ( .A(n2306), .Y(n2250) );
  CLKBUFX3 U405 ( .A(n2306), .Y(n2251) );
  CLKBUFX3 U406 ( .A(n2305), .Y(n2252) );
  CLKBUFX3 U407 ( .A(n2305), .Y(n2253) );
  CLKBUFX3 U408 ( .A(n2304), .Y(n2254) );
  CLKBUFX3 U409 ( .A(n2304), .Y(n2255) );
  CLKBUFX3 U410 ( .A(n2303), .Y(n2256) );
  CLKBUFX3 U411 ( .A(n2303), .Y(n2257) );
  CLKBUFX3 U412 ( .A(n2302), .Y(n2258) );
  CLKBUFX3 U413 ( .A(n2302), .Y(n2259) );
  CLKBUFX3 U414 ( .A(n2301), .Y(n2260) );
  CLKBUFX3 U415 ( .A(n2301), .Y(n2261) );
  CLKBUFX3 U416 ( .A(n2300), .Y(n2262) );
  CLKBUFX3 U417 ( .A(n2300), .Y(n2263) );
  CLKBUFX3 U418 ( .A(n2299), .Y(n2264) );
  CLKBUFX3 U419 ( .A(n2299), .Y(n2265) );
  CLKBUFX3 U420 ( .A(n2298), .Y(n2266) );
  CLKBUFX3 U421 ( .A(n2298), .Y(n2267) );
  CLKBUFX3 U422 ( .A(n2297), .Y(n2268) );
  CLKBUFX3 U423 ( .A(n2297), .Y(n2269) );
  CLKBUFX3 U424 ( .A(n2296), .Y(n2270) );
  CLKBUFX3 U425 ( .A(n2296), .Y(n2271) );
  CLKBUFX3 U426 ( .A(n2295), .Y(n2272) );
  CLKBUFX3 U427 ( .A(n2295), .Y(n2273) );
  CLKBUFX3 U428 ( .A(n2294), .Y(n2274) );
  CLKBUFX3 U429 ( .A(n2294), .Y(n2275) );
  CLKBUFX3 U430 ( .A(n2293), .Y(n2276) );
  CLKBUFX3 U431 ( .A(n2293), .Y(n2277) );
  CLKBUFX3 U432 ( .A(n2292), .Y(n2278) );
  CLKBUFX3 U433 ( .A(n2292), .Y(n2279) );
  CLKBUFX3 U434 ( .A(n2291), .Y(n2280) );
  CLKBUFX3 U435 ( .A(n2291), .Y(n2281) );
  CLKBUFX3 U436 ( .A(n2290), .Y(n2282) );
  CLKBUFX3 U437 ( .A(n2290), .Y(n2283) );
  CLKBUFX3 U438 ( .A(n2289), .Y(n2284) );
  CLKBUFX3 U439 ( .A(n2289), .Y(n2285) );
  CLKBUFX3 U440 ( .A(n2326), .Y(n2210) );
  CLKBUFX3 U441 ( .A(n2326), .Y(n2211) );
  CLKBUFX3 U442 ( .A(n2325), .Y(n2212) );
  CLKBUFX3 U443 ( .A(n2325), .Y(n2213) );
  CLKBUFX3 U444 ( .A(n2324), .Y(n2214) );
  CLKBUFX3 U445 ( .A(n2324), .Y(n2215) );
  CLKBUFX3 U446 ( .A(n2323), .Y(n2216) );
  CLKBUFX3 U447 ( .A(n2323), .Y(n2217) );
  CLKBUFX3 U448 ( .A(n2322), .Y(n2218) );
  CLKBUFX3 U449 ( .A(n2322), .Y(n2219) );
  CLKBUFX3 U450 ( .A(n2288), .Y(n2286) );
  CLKBUFX3 U451 ( .A(n2288), .Y(n2287) );
  CLKBUFX3 U452 ( .A(n471), .Y(n478) );
  CLKBUFX3 U453 ( .A(n469), .Y(n482) );
  CLKBUFX3 U454 ( .A(n467), .Y(n486) );
  CLKBUFX3 U455 ( .A(n465), .Y(n490) );
  CLKBUFX3 U456 ( .A(n463), .Y(n494) );
  CLKBUFX3 U457 ( .A(n470), .Y(n481) );
  CLKBUFX3 U458 ( .A(n469), .Y(n483) );
  CLKBUFX3 U459 ( .A(n468), .Y(n484) );
  CLKBUFX3 U460 ( .A(n468), .Y(n485) );
  CLKBUFX3 U461 ( .A(n467), .Y(n487) );
  CLKBUFX3 U462 ( .A(n466), .Y(n488) );
  CLKBUFX3 U463 ( .A(n466), .Y(n489) );
  CLKBUFX3 U464 ( .A(n465), .Y(n491) );
  CLKBUFX3 U465 ( .A(n464), .Y(n492) );
  CLKBUFX3 U466 ( .A(n464), .Y(n493) );
  CLKBUFX3 U467 ( .A(n472), .Y(n477) );
  CLKBUFX3 U468 ( .A(n472), .Y(n476) );
  CLKBUFX3 U469 ( .A(n463), .Y(n495) );
  CLKBUFX3 U470 ( .A(n471), .Y(n479) );
  CLKBUFX3 U471 ( .A(n470), .Y(n480) );
  CLKBUFX3 U472 ( .A(n899), .Y(n903) );
  CLKBUFX3 U473 ( .A(n899), .Y(n904) );
  CLKBUFX3 U474 ( .A(n898), .Y(n905) );
  CLKBUFX3 U475 ( .A(n898), .Y(n906) );
  CLKBUFX3 U476 ( .A(n897), .Y(n908) );
  CLKBUFX3 U477 ( .A(n897), .Y(n909) );
  CLKBUFX3 U478 ( .A(n896), .Y(n910) );
  CLKBUFX3 U479 ( .A(n896), .Y(n911) );
  CLKBUFX3 U480 ( .A(n895), .Y(n912) );
  CLKBUFX3 U481 ( .A(n895), .Y(n913) );
  CLKBUFX3 U482 ( .A(n894), .Y(n914) );
  CLKBUFX3 U483 ( .A(n894), .Y(n915) );
  CLKBUFX3 U484 ( .A(n893), .Y(n916) );
  CLKBUFX3 U485 ( .A(n893), .Y(n917) );
  CLKBUFX3 U486 ( .A(n892), .Y(n918) );
  CLKBUFX3 U487 ( .A(n892), .Y(n919) );
  CLKBUFX3 U488 ( .A(n891), .Y(n920) );
  CLKBUFX3 U489 ( .A(n891), .Y(n921) );
  CLKBUFX3 U490 ( .A(n890), .Y(n922) );
  CLKBUFX3 U491 ( .A(n890), .Y(n923) );
  CLKBUFX3 U492 ( .A(n2330), .Y(n2321) );
  CLKBUFX3 U493 ( .A(n2330), .Y(n2320) );
  CLKBUFX3 U494 ( .A(n2330), .Y(n2319) );
  CLKBUFX3 U495 ( .A(n2331), .Y(n2318) );
  CLKBUFX3 U496 ( .A(n2331), .Y(n2317) );
  CLKBUFX3 U497 ( .A(n2331), .Y(n2316) );
  CLKBUFX3 U498 ( .A(n2332), .Y(n2315) );
  CLKBUFX3 U499 ( .A(n2332), .Y(n2314) );
  CLKBUFX3 U500 ( .A(n2332), .Y(n2313) );
  CLKBUFX3 U501 ( .A(n2333), .Y(n2312) );
  CLKBUFX3 U502 ( .A(n2333), .Y(n2311) );
  CLKBUFX3 U503 ( .A(n2333), .Y(n2310) );
  CLKBUFX3 U504 ( .A(n2334), .Y(n2309) );
  CLKBUFX3 U505 ( .A(n2334), .Y(n2308) );
  CLKBUFX3 U506 ( .A(n2334), .Y(n2307) );
  CLKBUFX3 U507 ( .A(n2335), .Y(n2306) );
  CLKBUFX3 U508 ( .A(n2335), .Y(n2305) );
  CLKBUFX3 U509 ( .A(n2335), .Y(n2304) );
  CLKBUFX3 U510 ( .A(n2336), .Y(n2303) );
  CLKBUFX3 U511 ( .A(n2336), .Y(n2302) );
  CLKBUFX3 U512 ( .A(n2336), .Y(n2301) );
  CLKBUFX3 U513 ( .A(n2337), .Y(n2300) );
  CLKBUFX3 U514 ( .A(n2337), .Y(n2299) );
  CLKBUFX3 U515 ( .A(n2337), .Y(n2298) );
  CLKBUFX3 U516 ( .A(n2338), .Y(n2297) );
  CLKBUFX3 U517 ( .A(n2338), .Y(n2296) );
  CLKBUFX3 U518 ( .A(n2338), .Y(n2295) );
  CLKBUFX3 U519 ( .A(n2339), .Y(n2294) );
  CLKBUFX3 U520 ( .A(n2339), .Y(n2293) );
  CLKBUFX3 U521 ( .A(n2339), .Y(n2292) );
  CLKBUFX3 U522 ( .A(n2340), .Y(n2291) );
  CLKBUFX3 U523 ( .A(n2340), .Y(n2290) );
  CLKBUFX3 U524 ( .A(n2340), .Y(n2289) );
  CLKBUFX3 U525 ( .A(n430), .Y(n437) );
  CLKBUFX3 U526 ( .A(n428), .Y(n441) );
  CLKBUFX3 U527 ( .A(n426), .Y(n445) );
  CLKBUFX3 U528 ( .A(n424), .Y(n449) );
  CLKBUFX3 U529 ( .A(n422), .Y(n453) );
  CLKBUFX3 U530 ( .A(n429), .Y(n440) );
  CLKBUFX3 U531 ( .A(n428), .Y(n442) );
  CLKBUFX3 U532 ( .A(n427), .Y(n443) );
  CLKBUFX3 U533 ( .A(n427), .Y(n444) );
  CLKBUFX3 U534 ( .A(n426), .Y(n446) );
  CLKBUFX3 U535 ( .A(n425), .Y(n447) );
  CLKBUFX3 U536 ( .A(n425), .Y(n448) );
  CLKBUFX3 U537 ( .A(n424), .Y(n450) );
  CLKBUFX3 U538 ( .A(n423), .Y(n451) );
  CLKBUFX3 U539 ( .A(n423), .Y(n452) );
  CLKBUFX3 U540 ( .A(n431), .Y(n436) );
  CLKBUFX3 U541 ( .A(n431), .Y(n435) );
  CLKBUFX3 U542 ( .A(n422), .Y(n454) );
  CLKBUFX3 U543 ( .A(n430), .Y(n438) );
  CLKBUFX3 U544 ( .A(n429), .Y(n439) );
  CLKBUFX3 U545 ( .A(n856), .Y(n860) );
  CLKBUFX3 U546 ( .A(n856), .Y(n861) );
  CLKBUFX3 U547 ( .A(n855), .Y(n862) );
  CLKBUFX3 U548 ( .A(n855), .Y(n863) );
  CLKBUFX3 U549 ( .A(n854), .Y(n864) );
  CLKBUFX3 U550 ( .A(n854), .Y(n865) );
  CLKBUFX3 U551 ( .A(n853), .Y(n866) );
  CLKBUFX3 U552 ( .A(n853), .Y(n867) );
  CLKBUFX3 U553 ( .A(n852), .Y(n868) );
  CLKBUFX3 U554 ( .A(n852), .Y(n869) );
  CLKBUFX3 U555 ( .A(n851), .Y(n870) );
  CLKBUFX3 U556 ( .A(n851), .Y(n871) );
  CLKBUFX3 U557 ( .A(n850), .Y(n874) );
  CLKBUFX3 U558 ( .A(n850), .Y(n875) );
  CLKBUFX3 U559 ( .A(n849), .Y(n876) );
  CLKBUFX3 U560 ( .A(n849), .Y(n877) );
  CLKBUFX3 U561 ( .A(n848), .Y(n878) );
  CLKBUFX3 U562 ( .A(n848), .Y(n879) );
  CLKBUFX3 U563 ( .A(n847), .Y(n880) );
  CLKBUFX3 U564 ( .A(n847), .Y(n881) );
  CLKBUFX3 U565 ( .A(n2327), .Y(n2209) );
  CLKBUFX3 U566 ( .A(n2328), .Y(n2327) );
  CLKBUFX3 U567 ( .A(n473), .Y(n475) );
  CLKBUFX3 U568 ( .A(n900), .Y(n902) );
  CLKBUFX3 U569 ( .A(n1), .Y(n1024) );
  CLKBUFX3 U570 ( .A(n1), .Y(n1023) );
  CLKBUFX3 U571 ( .A(n2), .Y(n1019) );
  CLKBUFX3 U572 ( .A(n2), .Y(n1018) );
  CLKBUFX3 U573 ( .A(n3), .Y(n1016) );
  CLKBUFX3 U574 ( .A(n3), .Y(n1015) );
  CLKBUFX3 U575 ( .A(n6), .Y(n1013) );
  CLKBUFX3 U576 ( .A(n6), .Y(n1012) );
  CLKBUFX3 U577 ( .A(n8), .Y(n1010) );
  CLKBUFX3 U578 ( .A(n8), .Y(n1009) );
  CLKBUFX3 U579 ( .A(n10), .Y(n1007) );
  CLKBUFX3 U580 ( .A(n10), .Y(n1006) );
  CLKBUFX3 U581 ( .A(n12), .Y(n1004) );
  CLKBUFX3 U582 ( .A(n12), .Y(n1003) );
  CLKBUFX3 U583 ( .A(n14), .Y(n1001) );
  CLKBUFX3 U584 ( .A(n14), .Y(n1000) );
  CLKBUFX3 U585 ( .A(n16), .Y(n998) );
  CLKBUFX3 U586 ( .A(n16), .Y(n997) );
  CLKBUFX3 U587 ( .A(n18), .Y(n995) );
  CLKBUFX3 U588 ( .A(n18), .Y(n994) );
  CLKBUFX3 U589 ( .A(n20), .Y(n992) );
  CLKBUFX3 U590 ( .A(n20), .Y(n991) );
  CLKBUFX3 U591 ( .A(n22), .Y(n989) );
  CLKBUFX3 U592 ( .A(n22), .Y(n988) );
  CLKBUFX3 U593 ( .A(n24), .Y(n986) );
  CLKBUFX3 U594 ( .A(n24), .Y(n985) );
  CLKBUFX3 U595 ( .A(n26), .Y(n983) );
  CLKBUFX3 U596 ( .A(n26), .Y(n982) );
  CLKBUFX3 U597 ( .A(n28), .Y(n980) );
  CLKBUFX3 U598 ( .A(n28), .Y(n979) );
  CLKBUFX3 U599 ( .A(n30), .Y(n977) );
  CLKBUFX3 U600 ( .A(n30), .Y(n976) );
  CLKBUFX3 U601 ( .A(n32), .Y(n973) );
  CLKBUFX3 U602 ( .A(n32), .Y(n972) );
  CLKBUFX3 U603 ( .A(n34), .Y(n970) );
  CLKBUFX3 U604 ( .A(n34), .Y(n969) );
  CLKBUFX3 U605 ( .A(n36), .Y(n967) );
  CLKBUFX3 U606 ( .A(n36), .Y(n966) );
  CLKBUFX3 U607 ( .A(n38), .Y(n964) );
  CLKBUFX3 U608 ( .A(n38), .Y(n963) );
  CLKBUFX3 U609 ( .A(n40), .Y(n961) );
  CLKBUFX3 U610 ( .A(n40), .Y(n960) );
  CLKBUFX3 U611 ( .A(n42), .Y(n958) );
  CLKBUFX3 U612 ( .A(n42), .Y(n957) );
  CLKBUFX3 U613 ( .A(n44), .Y(n955) );
  CLKBUFX3 U614 ( .A(n44), .Y(n954) );
  CLKBUFX3 U615 ( .A(n46), .Y(n952) );
  CLKBUFX3 U616 ( .A(n46), .Y(n951) );
  CLKBUFX3 U617 ( .A(n48), .Y(n949) );
  CLKBUFX3 U618 ( .A(n48), .Y(n948) );
  CLKBUFX3 U619 ( .A(n50), .Y(n946) );
  CLKBUFX3 U620 ( .A(n50), .Y(n945) );
  CLKBUFX3 U621 ( .A(n52), .Y(n943) );
  CLKBUFX3 U622 ( .A(n52), .Y(n942) );
  CLKBUFX3 U623 ( .A(n54), .Y(n939) );
  CLKBUFX3 U624 ( .A(n54), .Y(n938) );
  CLKBUFX3 U625 ( .A(n56), .Y(n936) );
  CLKBUFX3 U626 ( .A(n56), .Y(n935) );
  CLKBUFX3 U627 ( .A(n58), .Y(n933) );
  CLKBUFX3 U628 ( .A(n58), .Y(n932) );
  CLKBUFX3 U629 ( .A(n60), .Y(n930) );
  CLKBUFX3 U630 ( .A(n60), .Y(n929) );
  CLKBUFX3 U631 ( .A(n62), .Y(n927) );
  CLKBUFX3 U632 ( .A(n62), .Y(n926) );
  CLKBUFX3 U633 ( .A(n2328), .Y(n2326) );
  CLKBUFX3 U634 ( .A(n2328), .Y(n2325) );
  CLKBUFX3 U635 ( .A(n2329), .Y(n2324) );
  CLKBUFX3 U636 ( .A(n2329), .Y(n2323) );
  CLKBUFX3 U637 ( .A(n2329), .Y(n2322) );
  CLKBUFX3 U638 ( .A(n2341), .Y(n2288) );
  CLKBUFX3 U639 ( .A(n2342), .Y(n2341) );
  CLKBUFX3 U640 ( .A(n1), .Y(n1025) );
  CLKBUFX3 U641 ( .A(n2), .Y(n1020) );
  CLKBUFX3 U642 ( .A(n3), .Y(n1017) );
  CLKBUFX3 U643 ( .A(n6), .Y(n1014) );
  CLKBUFX3 U644 ( .A(n8), .Y(n1011) );
  CLKBUFX3 U645 ( .A(n10), .Y(n1008) );
  CLKBUFX3 U646 ( .A(n12), .Y(n1005) );
  CLKBUFX3 U647 ( .A(n14), .Y(n1002) );
  CLKBUFX3 U648 ( .A(n16), .Y(n999) );
  CLKBUFX3 U649 ( .A(n18), .Y(n996) );
  CLKBUFX3 U650 ( .A(n20), .Y(n993) );
  CLKBUFX3 U651 ( .A(n22), .Y(n990) );
  CLKBUFX3 U652 ( .A(n24), .Y(n987) );
  CLKBUFX3 U653 ( .A(n26), .Y(n984) );
  CLKBUFX3 U654 ( .A(n28), .Y(n981) );
  CLKBUFX3 U655 ( .A(n30), .Y(n978) );
  CLKBUFX3 U656 ( .A(n32), .Y(n974) );
  CLKBUFX3 U657 ( .A(n34), .Y(n971) );
  CLKBUFX3 U658 ( .A(n36), .Y(n968) );
  CLKBUFX3 U659 ( .A(n38), .Y(n965) );
  CLKBUFX3 U660 ( .A(n40), .Y(n962) );
  CLKBUFX3 U661 ( .A(n42), .Y(n959) );
  CLKBUFX3 U662 ( .A(n44), .Y(n956) );
  CLKBUFX3 U663 ( .A(n46), .Y(n953) );
  CLKBUFX3 U664 ( .A(n48), .Y(n950) );
  CLKBUFX3 U665 ( .A(n50), .Y(n947) );
  CLKBUFX3 U666 ( .A(n52), .Y(n944) );
  CLKBUFX3 U667 ( .A(n54), .Y(n940) );
  CLKBUFX3 U668 ( .A(n56), .Y(n937) );
  CLKBUFX3 U669 ( .A(n58), .Y(n934) );
  CLKBUFX3 U670 ( .A(n60), .Y(n931) );
  CLKBUFX3 U671 ( .A(n62), .Y(n928) );
  CLKBUFX3 U672 ( .A(n458), .Y(n471) );
  CLKBUFX3 U673 ( .A(n417), .Y(n430) );
  CLKBUFX3 U674 ( .A(n459), .Y(n469) );
  CLKBUFX3 U675 ( .A(n418), .Y(n428) );
  CLKBUFX3 U676 ( .A(n460), .Y(n467) );
  CLKBUFX3 U677 ( .A(n419), .Y(n426) );
  CLKBUFX3 U678 ( .A(n461), .Y(n465) );
  CLKBUFX3 U679 ( .A(n420), .Y(n424) );
  CLKBUFX3 U680 ( .A(n462), .Y(n463) );
  CLKBUFX3 U681 ( .A(n421), .Y(n422) );
  CLKBUFX3 U682 ( .A(n459), .Y(n470) );
  CLKBUFX3 U683 ( .A(n418), .Y(n429) );
  CLKBUFX3 U684 ( .A(n460), .Y(n468) );
  CLKBUFX3 U685 ( .A(n419), .Y(n427) );
  CLKBUFX3 U686 ( .A(n461), .Y(n466) );
  CLKBUFX3 U687 ( .A(n420), .Y(n425) );
  CLKBUFX3 U688 ( .A(n462), .Y(n464) );
  CLKBUFX3 U689 ( .A(n421), .Y(n423) );
  CLKBUFX3 U690 ( .A(n458), .Y(n472) );
  CLKBUFX3 U691 ( .A(n417), .Y(n431) );
  CLKBUFX3 U692 ( .A(n885), .Y(n899) );
  CLKBUFX3 U693 ( .A(n842), .Y(n856) );
  CLKBUFX3 U694 ( .A(n885), .Y(n898) );
  CLKBUFX3 U695 ( .A(n842), .Y(n855) );
  CLKBUFX3 U696 ( .A(n886), .Y(n897) );
  CLKBUFX3 U697 ( .A(n843), .Y(n854) );
  CLKBUFX3 U698 ( .A(n886), .Y(n896) );
  CLKBUFX3 U699 ( .A(n843), .Y(n853) );
  CLKBUFX3 U700 ( .A(n887), .Y(n895) );
  CLKBUFX3 U701 ( .A(n844), .Y(n852) );
  CLKBUFX3 U702 ( .A(n887), .Y(n894) );
  CLKBUFX3 U703 ( .A(n844), .Y(n851) );
  CLKBUFX3 U704 ( .A(n888), .Y(n893) );
  CLKBUFX3 U705 ( .A(n845), .Y(n850) );
  CLKBUFX3 U706 ( .A(n888), .Y(n892) );
  CLKBUFX3 U707 ( .A(n845), .Y(n849) );
  CLKBUFX3 U708 ( .A(n889), .Y(n891) );
  CLKBUFX3 U709 ( .A(n846), .Y(n848) );
  CLKBUFX3 U710 ( .A(n889), .Y(n890) );
  CLKBUFX3 U711 ( .A(n846), .Y(n847) );
  CLKBUFX3 U712 ( .A(n432), .Y(n434) );
  CLKBUFX3 U713 ( .A(n857), .Y(n859) );
  CLKBUFX3 U714 ( .A(n2345), .Y(n2330) );
  CLKBUFX3 U715 ( .A(n2345), .Y(n2331) );
  CLKBUFX3 U716 ( .A(n2345), .Y(n2332) );
  CLKBUFX3 U717 ( .A(n2344), .Y(n2333) );
  CLKBUFX3 U718 ( .A(n2344), .Y(n2334) );
  CLKBUFX3 U719 ( .A(n2344), .Y(n2335) );
  CLKBUFX3 U720 ( .A(n2343), .Y(n2336) );
  CLKBUFX3 U721 ( .A(n2343), .Y(n2337) );
  CLKBUFX3 U722 ( .A(n2343), .Y(n2338) );
  CLKBUFX3 U723 ( .A(n2342), .Y(n2339) );
  CLKBUFX3 U724 ( .A(n2342), .Y(n2340) );
  CLKBUFX3 U725 ( .A(n473), .Y(n474) );
  CLKBUFX3 U726 ( .A(n900), .Y(n901) );
  CLKBUFX3 U727 ( .A(n432), .Y(n433) );
  CLKBUFX3 U728 ( .A(n857), .Y(n858) );
  CLKBUFX3 U729 ( .A(n1029), .Y(n1027) );
  CLKBUFX3 U730 ( .A(n1034), .Y(n1032) );
  CLKBUFX3 U731 ( .A(n1039), .Y(n1037) );
  CLKBUFX3 U732 ( .A(n2068), .Y(n1042) );
  CLKBUFX3 U733 ( .A(n2073), .Y(n2071) );
  CLKBUFX3 U734 ( .A(n2078), .Y(n2076) );
  CLKBUFX3 U735 ( .A(n2083), .Y(n2081) );
  CLKBUFX3 U736 ( .A(n2088), .Y(n2086) );
  CLKBUFX3 U737 ( .A(n2093), .Y(n2091) );
  CLKBUFX3 U738 ( .A(n2098), .Y(n2096) );
  CLKBUFX3 U739 ( .A(n2103), .Y(n2101) );
  CLKBUFX3 U740 ( .A(n2108), .Y(n2106) );
  CLKBUFX3 U741 ( .A(n2113), .Y(n2111) );
  CLKBUFX3 U742 ( .A(n2118), .Y(n2116) );
  CLKBUFX3 U743 ( .A(n2123), .Y(n2121) );
  CLKBUFX3 U744 ( .A(n2128), .Y(n2126) );
  CLKBUFX3 U745 ( .A(n2133), .Y(n2131) );
  CLKBUFX3 U746 ( .A(n2138), .Y(n2136) );
  CLKBUFX3 U747 ( .A(n2143), .Y(n2141) );
  CLKBUFX3 U748 ( .A(n2148), .Y(n2146) );
  CLKBUFX3 U749 ( .A(n2153), .Y(n2151) );
  CLKBUFX3 U750 ( .A(n2158), .Y(n2156) );
  CLKBUFX3 U751 ( .A(n2163), .Y(n2161) );
  CLKBUFX3 U752 ( .A(n1029), .Y(n1028) );
  CLKBUFX3 U753 ( .A(n1034), .Y(n1033) );
  CLKBUFX3 U754 ( .A(n1039), .Y(n1038) );
  CLKBUFX3 U755 ( .A(n2068), .Y(n1043) );
  CLKBUFX3 U756 ( .A(n2073), .Y(n2072) );
  CLKBUFX3 U757 ( .A(n2078), .Y(n2077) );
  CLKBUFX3 U758 ( .A(n2083), .Y(n2082) );
  CLKBUFX3 U759 ( .A(n2088), .Y(n2087) );
  CLKBUFX3 U760 ( .A(n2093), .Y(n2092) );
  CLKBUFX3 U761 ( .A(n2098), .Y(n2097) );
  CLKBUFX3 U762 ( .A(n2103), .Y(n2102) );
  CLKBUFX3 U763 ( .A(n2108), .Y(n2107) );
  CLKBUFX3 U764 ( .A(n2113), .Y(n2112) );
  CLKBUFX3 U765 ( .A(n2118), .Y(n2117) );
  CLKBUFX3 U766 ( .A(n2123), .Y(n2122) );
  CLKBUFX3 U767 ( .A(n2128), .Y(n2127) );
  CLKBUFX3 U768 ( .A(n2133), .Y(n2132) );
  CLKBUFX3 U769 ( .A(n2138), .Y(n2137) );
  CLKBUFX3 U770 ( .A(n2143), .Y(n2142) );
  CLKBUFX3 U771 ( .A(n2148), .Y(n2147) );
  CLKBUFX3 U772 ( .A(n2153), .Y(n2152) );
  CLKBUFX3 U773 ( .A(n2158), .Y(n2157) );
  CLKBUFX3 U774 ( .A(n2163), .Y(n2162) );
  NOR2BX1 U775 ( .AN(n7), .B(n1021), .Y(n6) );
  AND2X2 U776 ( .A(n872), .B(n206), .Y(n7) );
  NOR2BX1 U777 ( .AN(n9), .B(n1021), .Y(n8) );
  AND2X2 U778 ( .A(n872), .B(n172), .Y(n9) );
  NOR2BX1 U779 ( .AN(n11), .B(n1021), .Y(n10) );
  AND2X2 U780 ( .A(n872), .B(n138), .Y(n11) );
  NOR2BX1 U781 ( .AN(n13), .B(n1021), .Y(n12) );
  AND2X2 U782 ( .A(n872), .B(n104), .Y(n13) );
  NOR2BX1 U783 ( .AN(n15), .B(n1021), .Y(n14) );
  AND2X2 U784 ( .A(n872), .B(n70), .Y(n15) );
  NOR2BX1 U785 ( .AN(n17), .B(n1021), .Y(n16) );
  AND2X2 U786 ( .A(n607), .B(n308), .Y(n17) );
  NOR2BX1 U787 ( .AN(n19), .B(n1021), .Y(n18) );
  AND2X2 U788 ( .A(n607), .B(n274), .Y(n19) );
  NOR2BX1 U789 ( .AN(n21), .B(n1021), .Y(n20) );
  AND2X2 U790 ( .A(n607), .B(n240), .Y(n21) );
  NOR2BX1 U791 ( .AN(n23), .B(n1021), .Y(n22) );
  AND2X2 U792 ( .A(n607), .B(n206), .Y(n23) );
  NOR2BX1 U793 ( .AN(n25), .B(n1021), .Y(n24) );
  AND2X2 U794 ( .A(n607), .B(n172), .Y(n25) );
  NOR2BX1 U795 ( .AN(n27), .B(n1021), .Y(n26) );
  AND2X2 U796 ( .A(n607), .B(n138), .Y(n27) );
  NOR2BX1 U797 ( .AN(n29), .B(n1021), .Y(n28) );
  AND2X2 U798 ( .A(n607), .B(n104), .Y(n29) );
  NOR2BX1 U799 ( .AN(n31), .B(n1021), .Y(n30) );
  AND2X2 U800 ( .A(n607), .B(n70), .Y(n31) );
  NOR2BX1 U801 ( .AN(n33), .B(n1022), .Y(n32) );
  AND2X2 U802 ( .A(n342), .B(n308), .Y(n33) );
  NOR2BX1 U803 ( .AN(n35), .B(n1022), .Y(n34) );
  AND2X2 U804 ( .A(n342), .B(n274), .Y(n35) );
  NOR2BX1 U805 ( .AN(n37), .B(n1022), .Y(n36) );
  AND2X2 U806 ( .A(n342), .B(n240), .Y(n37) );
  NOR2BX1 U807 ( .AN(n39), .B(n1022), .Y(n38) );
  AND2X2 U808 ( .A(n342), .B(n206), .Y(n39) );
  NOR2BX1 U809 ( .AN(n41), .B(n1022), .Y(n40) );
  AND2X2 U810 ( .A(n342), .B(n172), .Y(n41) );
  NOR2BX1 U811 ( .AN(n43), .B(n1022), .Y(n42) );
  AND2X2 U812 ( .A(n342), .B(n138), .Y(n43) );
  NOR2BX1 U813 ( .AN(n45), .B(n1022), .Y(n44) );
  AND2X2 U814 ( .A(n342), .B(n104), .Y(n45) );
  NOR2BX1 U815 ( .AN(n47), .B(n1022), .Y(n46) );
  AND2X2 U816 ( .A(n342), .B(n70), .Y(n47) );
  NOR2BX1 U817 ( .AN(n49), .B(n1022), .Y(n48) );
  AND2X2 U818 ( .A(n308), .B(n69), .Y(n49) );
  NOR2BX1 U819 ( .AN(n51), .B(n1022), .Y(n50) );
  AND2X2 U820 ( .A(n274), .B(n69), .Y(n51) );
  NOR2BX1 U821 ( .AN(n53), .B(n1022), .Y(n52) );
  AND2X2 U822 ( .A(n240), .B(n69), .Y(n53) );
  NOR2BX1 U823 ( .AN(n55), .B(n1022), .Y(n54) );
  AND2X2 U824 ( .A(n206), .B(n69), .Y(n55) );
  NOR2BX1 U825 ( .AN(n57), .B(n1022), .Y(n56) );
  AND2X2 U826 ( .A(n172), .B(n69), .Y(n57) );
  NOR2BX1 U827 ( .AN(n59), .B(n1022), .Y(n58) );
  AND2X2 U828 ( .A(n138), .B(n69), .Y(n59) );
  NOR2BX1 U829 ( .AN(n61), .B(n1022), .Y(n60) );
  AND2X2 U830 ( .A(n104), .B(n69), .Y(n61) );
  NOR2BX1 U831 ( .AN(n63), .B(n1022), .Y(n62) );
  AND2X2 U832 ( .A(n69), .B(n70), .Y(n63) );
  CLKINVX1 U833 ( .A(n308), .Y(n2350) );
  CLKINVX1 U834 ( .A(n274), .Y(n2348) );
  CLKINVX1 U835 ( .A(n240), .Y(n2347) );
  CLKBUFX3 U836 ( .A(n406), .Y(n402) );
  CLKBUFX3 U837 ( .A(n407), .Y(n403) );
  CLKBUFX3 U838 ( .A(n407), .Y(n404) );
  CLKBUFX3 U839 ( .A(n405), .Y(n400) );
  CLKBUFX3 U840 ( .A(n406), .Y(n401) );
  CLKBUFX3 U841 ( .A(n830), .Y(n825) );
  CLKBUFX3 U842 ( .A(n831), .Y(n826) );
  CLKBUFX3 U843 ( .A(n831), .Y(n827) );
  CLKBUFX3 U844 ( .A(n832), .Y(n828) );
  CLKBUFX3 U845 ( .A(n832), .Y(n829) );
  CLKINVX1 U846 ( .A(n872), .Y(n2351) );
  CLKBUFX3 U847 ( .A(n839), .Y(n834) );
  CLKBUFX3 U848 ( .A(n839), .Y(n835) );
  CLKBUFX3 U849 ( .A(n840), .Y(n836) );
  CLKBUFX3 U850 ( .A(n840), .Y(n837) );
  CLKBUFX3 U851 ( .A(n2349), .Y(n1021) );
  CLKBUFX3 U852 ( .A(n2349), .Y(n1022) );
  CLKBUFX3 U853 ( .A(n405), .Y(n399) );
  CLKBUFX3 U854 ( .A(n830), .Y(n824) );
  CLKBUFX3 U855 ( .A(n496), .Y(n458) );
  CLKBUFX3 U856 ( .A(n455), .Y(n417) );
  CLKBUFX3 U857 ( .A(n496), .Y(n459) );
  CLKBUFX3 U858 ( .A(n455), .Y(n418) );
  CLKBUFX3 U859 ( .A(n497), .Y(n460) );
  CLKBUFX3 U860 ( .A(n456), .Y(n419) );
  CLKBUFX3 U861 ( .A(n497), .Y(n461) );
  CLKBUFX3 U862 ( .A(n456), .Y(n420) );
  CLKBUFX3 U863 ( .A(n497), .Y(n462) );
  CLKBUFX3 U864 ( .A(n456), .Y(n421) );
  CLKBUFX3 U865 ( .A(n924), .Y(n885) );
  CLKBUFX3 U866 ( .A(n882), .Y(n842) );
  CLKBUFX3 U867 ( .A(n924), .Y(n886) );
  CLKBUFX3 U868 ( .A(n882), .Y(n843) );
  CLKBUFX3 U869 ( .A(n925), .Y(n887) );
  CLKBUFX3 U870 ( .A(n883), .Y(n844) );
  CLKBUFX3 U871 ( .A(n925), .Y(n888) );
  CLKBUFX3 U872 ( .A(n883), .Y(n845) );
  CLKBUFX3 U873 ( .A(n925), .Y(n889) );
  CLKBUFX3 U874 ( .A(n883), .Y(n846) );
  CLKBUFX3 U875 ( .A(n457), .Y(n473) );
  CLKBUFX3 U876 ( .A(n496), .Y(n457) );
  CLKBUFX3 U877 ( .A(n416), .Y(n432) );
  CLKBUFX3 U878 ( .A(n455), .Y(n416) );
  CLKBUFX3 U879 ( .A(n884), .Y(n900) );
  CLKBUFX3 U880 ( .A(n924), .Y(n884) );
  CLKBUFX3 U881 ( .A(n841), .Y(n857) );
  CLKBUFX3 U882 ( .A(n882), .Y(n841) );
  CLKBUFX3 U883 ( .A(n2207), .Y(n2345) );
  CLKBUFX3 U884 ( .A(n2207), .Y(n2344) );
  CLKBUFX3 U885 ( .A(n2206), .Y(n2343) );
  CLKBUFX3 U886 ( .A(n2206), .Y(n2342) );
  CLKBUFX3 U887 ( .A(n2346), .Y(n2328) );
  CLKBUFX3 U888 ( .A(n2346), .Y(n2329) );
  CLKBUFX3 U889 ( .A(WriteData_i[0]), .Y(n1029) );
  CLKBUFX3 U890 ( .A(WriteData_i[1]), .Y(n1034) );
  CLKBUFX3 U891 ( .A(WriteData_i[2]), .Y(n1039) );
  CLKBUFX3 U892 ( .A(WriteData_i[3]), .Y(n2068) );
  CLKBUFX3 U893 ( .A(WriteData_i[4]), .Y(n2073) );
  CLKBUFX3 U894 ( .A(WriteData_i[5]), .Y(n2078) );
  CLKBUFX3 U895 ( .A(WriteData_i[6]), .Y(n2083) );
  CLKBUFX3 U896 ( .A(WriteData_i[7]), .Y(n2088) );
  CLKBUFX3 U897 ( .A(WriteData_i[8]), .Y(n2093) );
  CLKBUFX3 U898 ( .A(WriteData_i[9]), .Y(n2098) );
  CLKBUFX3 U899 ( .A(WriteData_i[10]), .Y(n2103) );
  CLKBUFX3 U900 ( .A(WriteData_i[11]), .Y(n2108) );
  CLKBUFX3 U901 ( .A(WriteData_i[12]), .Y(n2113) );
  CLKBUFX3 U902 ( .A(WriteData_i[13]), .Y(n2118) );
  CLKBUFX3 U903 ( .A(WriteData_i[14]), .Y(n2123) );
  CLKBUFX3 U904 ( .A(WriteData_i[15]), .Y(n2128) );
  CLKBUFX3 U905 ( .A(WriteData_i[16]), .Y(n2133) );
  CLKBUFX3 U906 ( .A(WriteData_i[17]), .Y(n2138) );
  CLKBUFX3 U907 ( .A(WriteData_i[18]), .Y(n2143) );
  CLKBUFX3 U908 ( .A(WriteData_i[19]), .Y(n2148) );
  CLKBUFX3 U909 ( .A(WriteData_i[20]), .Y(n2153) );
  CLKBUFX3 U910 ( .A(WriteData_i[21]), .Y(n2158) );
  CLKBUFX3 U911 ( .A(WriteData_i[22]), .Y(n2163) );
  CLKBUFX3 U912 ( .A(WriteData_i[23]), .Y(n2168) );
  CLKBUFX3 U913 ( .A(WriteData_i[24]), .Y(n2173) );
  CLKBUFX3 U914 ( .A(WriteData_i[25]), .Y(n2178) );
  CLKBUFX3 U915 ( .A(WriteData_i[26]), .Y(n2183) );
  CLKBUFX3 U916 ( .A(WriteData_i[27]), .Y(n2188) );
  CLKBUFX3 U917 ( .A(WriteData_i[28]), .Y(n2193) );
  CLKBUFX3 U918 ( .A(WriteData_i[29]), .Y(n2198) );
  CLKBUFX3 U919 ( .A(WriteData_i[30]), .Y(n2203) );
  CLKBUFX3 U920 ( .A(n1030), .Y(n1026) );
  CLKBUFX3 U921 ( .A(WriteData_i[0]), .Y(n1030) );
  CLKBUFX3 U922 ( .A(n1035), .Y(n1031) );
  CLKBUFX3 U923 ( .A(WriteData_i[1]), .Y(n1035) );
  CLKBUFX3 U924 ( .A(n1040), .Y(n1036) );
  CLKBUFX3 U925 ( .A(WriteData_i[2]), .Y(n1040) );
  CLKBUFX3 U926 ( .A(n2069), .Y(n1041) );
  CLKBUFX3 U927 ( .A(WriteData_i[3]), .Y(n2069) );
  CLKBUFX3 U928 ( .A(n2074), .Y(n2070) );
  CLKBUFX3 U929 ( .A(WriteData_i[4]), .Y(n2074) );
  CLKBUFX3 U930 ( .A(n2079), .Y(n2075) );
  CLKBUFX3 U931 ( .A(WriteData_i[5]), .Y(n2079) );
  CLKBUFX3 U932 ( .A(n2084), .Y(n2080) );
  CLKBUFX3 U933 ( .A(WriteData_i[6]), .Y(n2084) );
  CLKBUFX3 U934 ( .A(n2089), .Y(n2085) );
  CLKBUFX3 U935 ( .A(WriteData_i[7]), .Y(n2089) );
  CLKBUFX3 U936 ( .A(n2094), .Y(n2090) );
  CLKBUFX3 U937 ( .A(WriteData_i[8]), .Y(n2094) );
  CLKBUFX3 U938 ( .A(n2099), .Y(n2095) );
  CLKBUFX3 U939 ( .A(WriteData_i[9]), .Y(n2099) );
  CLKBUFX3 U940 ( .A(n2104), .Y(n2100) );
  CLKBUFX3 U941 ( .A(WriteData_i[10]), .Y(n2104) );
  CLKBUFX3 U942 ( .A(n2109), .Y(n2105) );
  CLKBUFX3 U943 ( .A(WriteData_i[11]), .Y(n2109) );
  CLKBUFX3 U944 ( .A(n2114), .Y(n2110) );
  CLKBUFX3 U945 ( .A(WriteData_i[12]), .Y(n2114) );
  CLKBUFX3 U946 ( .A(n2119), .Y(n2115) );
  CLKBUFX3 U947 ( .A(WriteData_i[13]), .Y(n2119) );
  CLKBUFX3 U948 ( .A(n2124), .Y(n2120) );
  CLKBUFX3 U949 ( .A(WriteData_i[14]), .Y(n2124) );
  CLKBUFX3 U950 ( .A(n2129), .Y(n2125) );
  CLKBUFX3 U951 ( .A(WriteData_i[15]), .Y(n2129) );
  CLKBUFX3 U952 ( .A(n2134), .Y(n2130) );
  CLKBUFX3 U953 ( .A(WriteData_i[16]), .Y(n2134) );
  CLKBUFX3 U954 ( .A(n2139), .Y(n2135) );
  CLKBUFX3 U955 ( .A(WriteData_i[17]), .Y(n2139) );
  CLKBUFX3 U956 ( .A(n2144), .Y(n2140) );
  CLKBUFX3 U957 ( .A(WriteData_i[18]), .Y(n2144) );
  CLKBUFX3 U958 ( .A(n2149), .Y(n2145) );
  CLKBUFX3 U959 ( .A(WriteData_i[19]), .Y(n2149) );
  CLKBUFX3 U960 ( .A(n2154), .Y(n2150) );
  CLKBUFX3 U961 ( .A(WriteData_i[20]), .Y(n2154) );
  CLKBUFX3 U962 ( .A(n2159), .Y(n2155) );
  CLKBUFX3 U963 ( .A(WriteData_i[21]), .Y(n2159) );
  CLKBUFX3 U964 ( .A(n2164), .Y(n2160) );
  CLKBUFX3 U965 ( .A(WriteData_i[22]), .Y(n2164) );
  CLKBUFX3 U966 ( .A(n2169), .Y(n2165) );
  CLKBUFX3 U967 ( .A(WriteData_i[23]), .Y(n2169) );
  CLKBUFX3 U968 ( .A(n2174), .Y(n2170) );
  CLKBUFX3 U969 ( .A(WriteData_i[24]), .Y(n2174) );
  CLKBUFX3 U970 ( .A(n2179), .Y(n2175) );
  CLKBUFX3 U971 ( .A(WriteData_i[25]), .Y(n2179) );
  CLKBUFX3 U972 ( .A(n2184), .Y(n2180) );
  CLKBUFX3 U973 ( .A(WriteData_i[26]), .Y(n2184) );
  CLKBUFX3 U974 ( .A(n2189), .Y(n2185) );
  CLKBUFX3 U975 ( .A(WriteData_i[27]), .Y(n2189) );
  CLKBUFX3 U976 ( .A(n2194), .Y(n2190) );
  CLKBUFX3 U977 ( .A(WriteData_i[28]), .Y(n2194) );
  CLKBUFX3 U978 ( .A(n2199), .Y(n2195) );
  CLKBUFX3 U979 ( .A(WriteData_i[29]), .Y(n2199) );
  CLKBUFX3 U980 ( .A(n2204), .Y(n2200) );
  CLKBUFX3 U981 ( .A(WriteData_i[30]), .Y(n2204) );
  AND2X2 U982 ( .A(Reg_W_i[4]), .B(n2355), .Y(n607) );
  AND2X2 U983 ( .A(Reg_W_i[4]), .B(Reg_W_i[3]), .Y(n872) );
  AND2X2 U984 ( .A(Reg_W_i[2]), .B(n873), .Y(n206) );
  AND2X2 U985 ( .A(Reg_W_i[2]), .B(n975), .Y(n308) );
  AND2X2 U986 ( .A(Reg_W_i[2]), .B(n941), .Y(n274) );
  AND2X2 U987 ( .A(Reg_W_i[2]), .B(n907), .Y(n240) );
  CLKINVX1 U988 ( .A(RegWrite_i), .Y(n2349) );
  NOR2X1 U989 ( .A(n2354), .B(Reg_W_i[1]), .Y(n907) );
  NOR2X1 U990 ( .A(Reg_W_i[0]), .B(Reg_W_i[1]), .Y(n873) );
  CLKBUFX3 U991 ( .A(n398), .Y(n395) );
  CLKBUFX3 U992 ( .A(n398), .Y(n396) );
  CLKBUFX3 U993 ( .A(n823), .Y(n820) );
  CLKBUFX3 U994 ( .A(n823), .Y(n821) );
  CLKINVX1 U995 ( .A(Reg_W_i[0]), .Y(n2354) );
  CLKINVX1 U996 ( .A(Reg_W_i[3]), .Y(n2355) );
  CLKBUFX3 U997 ( .A(n414), .Y(n410) );
  CLKBUFX3 U998 ( .A(n415), .Y(n411) );
  CLKBUFX3 U999 ( .A(n415), .Y(n412) );
  CLKBUFX3 U1000 ( .A(n414), .Y(n409) );
  CLKBUFX3 U1001 ( .A(n838), .Y(n833) );
  CLKBUFX3 U1002 ( .A(N474), .Y(n838) );
  AND2X2 U1003 ( .A(Reg_W_i[1]), .B(Reg_W_i[0]), .Y(n975) );
  AND2X2 U1004 ( .A(Reg_W_i[1]), .B(n2354), .Y(n941) );
  CLKBUFX3 U1005 ( .A(rst_n), .Y(n2207) );
  CLKBUFX3 U1006 ( .A(rst_n), .Y(n2206) );
  CLKBUFX3 U1007 ( .A(N470), .Y(n405) );
  CLKBUFX3 U1008 ( .A(N470), .Y(n406) );
  CLKBUFX3 U1009 ( .A(N470), .Y(n407) );
  CLKBUFX3 U1010 ( .A(N475), .Y(n830) );
  CLKBUFX3 U1011 ( .A(N474), .Y(n839) );
  CLKBUFX3 U1012 ( .A(N475), .Y(n831) );
  CLKBUFX3 U1013 ( .A(N475), .Y(n832) );
  CLKBUFX3 U1014 ( .A(N474), .Y(n840) );
  CLKBUFX3 U1015 ( .A(N467), .Y(n496) );
  CLKBUFX3 U1016 ( .A(N468), .Y(n455) );
  CLKBUFX3 U1017 ( .A(N467), .Y(n497) );
  CLKBUFX3 U1018 ( .A(N468), .Y(n456) );
  CLKBUFX3 U1019 ( .A(N472), .Y(n924) );
  CLKBUFX3 U1020 ( .A(N473), .Y(n882) );
  CLKBUFX3 U1021 ( .A(N472), .Y(n925) );
  CLKBUFX3 U1022 ( .A(N473), .Y(n883) );
  CLKBUFX3 U1023 ( .A(n2208), .Y(n2346) );
  CLKBUFX3 U1024 ( .A(rst_n), .Y(n2208) );
  MX4X1 U1025 ( .A(n171), .B(n169), .C(n170), .D(n168), .S0(n400), .S1(n408), 
        .Y(n86) );
  MX4X1 U1026 ( .A(n167), .B(n165), .C(n166), .D(n164), .S0(n400), .S1(n408), 
        .Y(n87) );
  MX4X1 U1027 ( .A(n188), .B(n186), .C(n187), .D(n185), .S0(n400), .S1(n409), 
        .Y(n90) );
  MX4X1 U1028 ( .A(n184), .B(n182), .C(n183), .D(n181), .S0(n400), .S1(n409), 
        .Y(n91) );
  MX4X1 U1029 ( .A(n196), .B(n194), .C(n195), .D(n193), .S0(n400), .S1(n409), 
        .Y(n92) );
  MX4X1 U1030 ( .A(n192), .B(n190), .C(n191), .D(n189), .S0(n400), .S1(n409), 
        .Y(n93) );
  MXI4X1 U1031 ( .A(\register[0][7] ), .B(\register[1][7] ), .C(
        \register[2][7] ), .D(\register[3][7] ), .S0(n479), .S1(n438), .Y(n196) );
  MX4X1 U1032 ( .A(n155), .B(n153), .C(n154), .D(n152), .S0(n400), .S1(n408), 
        .Y(n82) );
  MX4X1 U1033 ( .A(n151), .B(n149), .C(n150), .D(n148), .S0(n400), .S1(n408), 
        .Y(n83) );
  MX4X1 U1034 ( .A(n180), .B(n178), .C(n179), .D(n177), .S0(n400), .S1(n408), 
        .Y(n88) );
  MX4X1 U1035 ( .A(n176), .B(n174), .C(n175), .D(n173), .S0(n400), .S1(n408), 
        .Y(n89) );
  MXI2X2 U1036 ( .A(n80), .B(n81), .S0(n394), .Y(ReadData1_o[0]) );
  MX4X1 U1037 ( .A(n139), .B(n136), .C(n137), .D(n135), .S0(n399), .S1(n408), 
        .Y(n80) );
  MX4X1 U1038 ( .A(n134), .B(n132), .C(n133), .D(n131), .S0(n399), .S1(n408), 
        .Y(n81) );
  MXI2X1 U1039 ( .A(n502), .B(n503), .S0(n819), .Y(ReadData2_o[2]) );
  MX4X1 U1040 ( .A(n581), .B(n579), .C(n580), .D(n578), .S0(n825), .S1(n833), 
        .Y(n503) );
  MX4X1 U1041 ( .A(n585), .B(n583), .C(n584), .D(n582), .S0(n825), .S1(n833), 
        .Y(n502) );
  MXI2X1 U1042 ( .A(n500), .B(n501), .S0(n819), .Y(ReadData2_o[1]) );
  MX4X1 U1043 ( .A(n573), .B(n571), .C(n572), .D(n570), .S0(n824), .S1(n833), 
        .Y(n501) );
  MXI2X1 U1044 ( .A(n498), .B(n499), .S0(n819), .Y(ReadData2_o[0]) );
  MX4X1 U1045 ( .A(n565), .B(n563), .C(n564), .D(n562), .S0(n824), .S1(n833), 
        .Y(n499) );
  MX4X1 U1046 ( .A(n589), .B(n587), .C(n588), .D(n586), .S0(n825), .S1(n833), 
        .Y(n505) );
  MX4X1 U1047 ( .A(n593), .B(n591), .C(n592), .D(n590), .S0(n825), .S1(n833), 
        .Y(n504) );
  MX4X1 U1048 ( .A(n597), .B(n595), .C(n596), .D(n594), .S0(n825), .S1(n833), 
        .Y(n507) );
  MX4X1 U1049 ( .A(n601), .B(n599), .C(n600), .D(n598), .S0(n825), .S1(n833), 
        .Y(n506) );
  MXI4X1 U1050 ( .A(\register[28][4] ), .B(\register[29][4] ), .C(
        \register[30][4] ), .D(\register[31][4] ), .S0(n904), .S1(n861), .Y(
        n594) );
  MX4X1 U1051 ( .A(n605), .B(n603), .C(n604), .D(n602), .S0(n825), .S1(n833), 
        .Y(n509) );
  MX4X1 U1052 ( .A(n610), .B(n608), .C(n609), .D(n606), .S0(n825), .S1(n833), 
        .Y(n508) );
  MXI4X1 U1053 ( .A(\register[28][5] ), .B(\register[29][5] ), .C(
        \register[30][5] ), .D(\register[31][5] ), .S0(n905), .S1(n862), .Y(
        n602) );
  MX4X1 U1054 ( .A(n614), .B(n612), .C(n613), .D(n611), .S0(n825), .S1(n834), 
        .Y(n511) );
  MX4X1 U1055 ( .A(n618), .B(n616), .C(n617), .D(n615), .S0(n825), .S1(n834), 
        .Y(n510) );
  MXI4X1 U1056 ( .A(\register[28][6] ), .B(\register[29][6] ), .C(
        \register[30][6] ), .D(\register[31][6] ), .S0(n905), .S1(n862), .Y(
        n611) );
  MXI2X1 U1057 ( .A(n512), .B(n513), .S0(n819), .Y(ReadData2_o[7]) );
  MX4X1 U1058 ( .A(n622), .B(n620), .C(n621), .D(n619), .S0(n825), .S1(n834), 
        .Y(n513) );
  MX4X1 U1059 ( .A(n626), .B(n624), .C(n625), .D(n623), .S0(n825), .S1(n834), 
        .Y(n512) );
  MXI4X1 U1060 ( .A(\register[28][7] ), .B(\register[29][7] ), .C(
        \register[30][7] ), .D(\register[31][7] ), .S0(n906), .S1(n863), .Y(
        n619) );
  MXI2X1 U1061 ( .A(n514), .B(n515), .S0(n820), .Y(ReadData2_o[8]) );
  MX4X1 U1062 ( .A(n630), .B(n628), .C(n629), .D(n627), .S0(n826), .S1(n834), 
        .Y(n515) );
  MX4X1 U1063 ( .A(n634), .B(n632), .C(n633), .D(n631), .S0(n826), .S1(n834), 
        .Y(n514) );
  MXI4X1 U1064 ( .A(\register[28][8] ), .B(\register[29][8] ), .C(
        \register[30][8] ), .D(\register[31][8] ), .S0(n908), .S1(n864), .Y(
        n627) );
  MX4X1 U1065 ( .A(n200), .B(n198), .C(n199), .D(n197), .S0(n401), .S1(n409), 
        .Y(n95) );
  MX4X1 U1066 ( .A(n204), .B(n202), .C(n203), .D(n201), .S0(n401), .S1(n409), 
        .Y(n94) );
  MXI4X1 U1067 ( .A(\register[28][8] ), .B(\register[29][8] ), .C(
        \register[30][8] ), .D(\register[31][8] ), .S0(n480), .S1(n439), .Y(
        n197) );
  MX4X1 U1068 ( .A(n163), .B(n161), .C(n162), .D(n160), .S0(n400), .S1(n408), 
        .Y(n84) );
  MX4X1 U1069 ( .A(n159), .B(n157), .C(n158), .D(n156), .S0(n400), .S1(n408), 
        .Y(n85) );
  MXI4X1 U1070 ( .A(\register[20][7] ), .B(\register[21][7] ), .C(
        \register[22][7] ), .D(\register[23][7] ), .S0(n479), .S1(n438), .Y(
        n191) );
  MXI4X1 U1071 ( .A(\register[4][7] ), .B(\register[5][7] ), .C(
        \register[6][7] ), .D(\register[7][7] ), .S0(n479), .S1(n438), .Y(n195) );
  MXI4X1 U1072 ( .A(\register[4][8] ), .B(\register[5][8] ), .C(
        \register[6][8] ), .D(\register[7][8] ), .S0(n480), .S1(n439), .Y(n203) );
  MXI4X1 U1073 ( .A(\register[20][8] ), .B(\register[21][8] ), .C(
        \register[22][8] ), .D(\register[23][8] ), .S0(n480), .S1(n439), .Y(
        n199) );
  MXI4X1 U1074 ( .A(\register[4][4] ), .B(\register[5][4] ), .C(
        \register[6][4] ), .D(\register[7][4] ), .S0(n904), .S1(n861), .Y(n600) );
  MXI4X1 U1075 ( .A(\register[20][4] ), .B(\register[21][4] ), .C(
        \register[22][4] ), .D(\register[23][4] ), .S0(n904), .S1(n861), .Y(
        n596) );
  MXI4X1 U1076 ( .A(\register[4][5] ), .B(\register[5][5] ), .C(
        \register[6][5] ), .D(\register[7][5] ), .S0(n905), .S1(n862), .Y(n609) );
  MXI4X1 U1077 ( .A(\register[20][5] ), .B(\register[21][5] ), .C(
        \register[22][5] ), .D(\register[23][5] ), .S0(n905), .S1(n862), .Y(
        n604) );
  MXI4X1 U1078 ( .A(\register[4][6] ), .B(\register[5][6] ), .C(
        \register[6][6] ), .D(\register[7][6] ), .S0(n906), .S1(n863), .Y(n617) );
  MXI4X1 U1079 ( .A(\register[20][6] ), .B(\register[21][6] ), .C(
        \register[22][6] ), .D(\register[23][6] ), .S0(n905), .S1(n862), .Y(
        n613) );
  MXI4X1 U1080 ( .A(\register[4][7] ), .B(\register[5][7] ), .C(
        \register[6][7] ), .D(\register[7][7] ), .S0(n906), .S1(n863), .Y(n625) );
  MXI4X1 U1081 ( .A(\register[20][7] ), .B(\register[21][7] ), .C(
        \register[22][7] ), .D(\register[23][7] ), .S0(n906), .S1(n863), .Y(
        n621) );
  MXI4X1 U1082 ( .A(\register[4][8] ), .B(\register[5][8] ), .C(
        \register[6][8] ), .D(\register[7][8] ), .S0(n908), .S1(n864), .Y(n633) );
  MXI4X1 U1083 ( .A(\register[20][8] ), .B(\register[21][8] ), .C(
        \register[22][8] ), .D(\register[23][8] ), .S0(n908), .S1(n864), .Y(
        n629) );
  MXI4X1 U1084 ( .A(\register[16][7] ), .B(\register[17][7] ), .C(
        \register[18][7] ), .D(\register[19][7] ), .S0(n479), .S1(n438), .Y(
        n192) );
  MXI4X1 U1085 ( .A(\register[0][8] ), .B(\register[1][8] ), .C(
        \register[2][8] ), .D(\register[3][8] ), .S0(n480), .S1(n439), .Y(n204) );
  MXI4X1 U1086 ( .A(\register[16][8] ), .B(\register[17][8] ), .C(
        \register[18][8] ), .D(\register[19][8] ), .S0(n480), .S1(n439), .Y(
        n200) );
  MXI4X1 U1087 ( .A(\register[0][4] ), .B(\register[1][4] ), .C(
        \register[2][4] ), .D(\register[3][4] ), .S0(n904), .S1(n861), .Y(n601) );
  MXI4X1 U1088 ( .A(\register[16][4] ), .B(\register[17][4] ), .C(
        \register[18][4] ), .D(\register[19][4] ), .S0(n904), .S1(n861), .Y(
        n597) );
  MXI4X1 U1089 ( .A(\register[0][5] ), .B(\register[1][5] ), .C(
        \register[2][5] ), .D(\register[3][5] ), .S0(n905), .S1(n862), .Y(n610) );
  MXI4X1 U1090 ( .A(\register[16][5] ), .B(\register[17][5] ), .C(
        \register[18][5] ), .D(\register[19][5] ), .S0(n905), .S1(n862), .Y(
        n605) );
  MXI4X1 U1091 ( .A(\register[0][6] ), .B(\register[1][6] ), .C(
        \register[2][6] ), .D(\register[3][6] ), .S0(n906), .S1(n863), .Y(n618) );
  MXI4X1 U1092 ( .A(\register[16][6] ), .B(\register[17][6] ), .C(
        \register[18][6] ), .D(\register[19][6] ), .S0(n905), .S1(n862), .Y(
        n614) );
  MXI4X1 U1093 ( .A(\register[0][7] ), .B(\register[1][7] ), .C(
        \register[2][7] ), .D(\register[3][7] ), .S0(n906), .S1(n863), .Y(n626) );
  MXI4X1 U1094 ( .A(\register[16][7] ), .B(\register[17][7] ), .C(
        \register[18][7] ), .D(\register[19][7] ), .S0(n906), .S1(n863), .Y(
        n622) );
  MXI4X1 U1095 ( .A(\register[0][8] ), .B(\register[1][8] ), .C(
        \register[2][8] ), .D(\register[3][8] ), .S0(n908), .S1(n864), .Y(n634) );
  MXI4X1 U1096 ( .A(\register[16][8] ), .B(\register[17][8] ), .C(
        \register[18][8] ), .D(\register[19][8] ), .S0(n908), .S1(n864), .Y(
        n630) );
  MX4X1 U1097 ( .A(n2353), .B(n2352), .C(n64), .D(n65), .S0(n474), .S1(n433), 
        .Y(n131) );
  MXI4X1 U1098 ( .A(\register[28][7] ), .B(\register[29][7] ), .C(
        \register[30][7] ), .D(\register[31][7] ), .S0(n479), .S1(n438), .Y(
        n189) );
  MXI4X1 U1099 ( .A(\register[12][7] ), .B(\register[13][7] ), .C(
        \register[14][7] ), .D(\register[15][7] ), .S0(n479), .S1(n438), .Y(
        n193) );
  MXI4X1 U1100 ( .A(\register[12][8] ), .B(\register[13][8] ), .C(
        \register[14][8] ), .D(\register[15][8] ), .S0(n480), .S1(n439), .Y(
        n201) );
  MXI4X1 U1101 ( .A(\register[12][4] ), .B(\register[13][4] ), .C(
        \register[14][4] ), .D(\register[15][4] ), .S0(n904), .S1(n861), .Y(
        n598) );
  MXI4X1 U1102 ( .A(\register[12][5] ), .B(\register[13][5] ), .C(
        \register[14][5] ), .D(\register[15][5] ), .S0(n905), .S1(n862), .Y(
        n606) );
  MXI4X1 U1103 ( .A(\register[12][6] ), .B(\register[13][6] ), .C(
        \register[14][6] ), .D(\register[15][6] ), .S0(n906), .S1(n863), .Y(
        n615) );
  MXI4X1 U1104 ( .A(\register[12][7] ), .B(\register[13][7] ), .C(
        \register[14][7] ), .D(\register[15][7] ), .S0(n906), .S1(n863), .Y(
        n623) );
  MXI4X1 U1105 ( .A(\register[12][8] ), .B(\register[13][8] ), .C(
        \register[14][8] ), .D(\register[15][8] ), .S0(n908), .S1(n864), .Y(
        n631) );
  MXI4X1 U1106 ( .A(\register[24][7] ), .B(\register[25][7] ), .C(
        \register[26][7] ), .D(\register[27][7] ), .S0(n479), .S1(n438), .Y(
        n190) );
  MXI4X1 U1107 ( .A(\register[8][7] ), .B(\register[9][7] ), .C(
        \register[10][7] ), .D(\register[11][7] ), .S0(n479), .S1(n438), .Y(
        n194) );
  MXI4X1 U1108 ( .A(\register[8][8] ), .B(\register[9][8] ), .C(
        \register[10][8] ), .D(\register[11][8] ), .S0(n480), .S1(n439), .Y(
        n202) );
  MXI4X1 U1109 ( .A(\register[24][8] ), .B(\register[25][8] ), .C(
        \register[26][8] ), .D(\register[27][8] ), .S0(n480), .S1(n439), .Y(
        n198) );
  MXI4X1 U1110 ( .A(\register[8][4] ), .B(\register[9][4] ), .C(
        \register[10][4] ), .D(\register[11][4] ), .S0(n904), .S1(n861), .Y(
        n599) );
  MXI4X1 U1111 ( .A(\register[24][4] ), .B(\register[25][4] ), .C(
        \register[26][4] ), .D(\register[27][4] ), .S0(n904), .S1(n861), .Y(
        n595) );
  MXI4X1 U1112 ( .A(\register[8][5] ), .B(\register[9][5] ), .C(
        \register[10][5] ), .D(\register[11][5] ), .S0(n905), .S1(n862), .Y(
        n608) );
  MXI4X1 U1113 ( .A(\register[24][5] ), .B(\register[25][5] ), .C(
        \register[26][5] ), .D(\register[27][5] ), .S0(n905), .S1(n862), .Y(
        n603) );
  MXI4X1 U1114 ( .A(\register[8][6] ), .B(\register[9][6] ), .C(
        \register[10][6] ), .D(\register[11][6] ), .S0(n906), .S1(n863), .Y(
        n616) );
  MXI4X1 U1115 ( .A(\register[24][6] ), .B(\register[25][6] ), .C(
        \register[26][6] ), .D(\register[27][6] ), .S0(n905), .S1(n862), .Y(
        n612) );
  MXI4X1 U1116 ( .A(\register[8][7] ), .B(\register[9][7] ), .C(
        \register[10][7] ), .D(\register[11][7] ), .S0(n906), .S1(n863), .Y(
        n624) );
  MXI4X1 U1117 ( .A(\register[24][7] ), .B(\register[25][7] ), .C(
        \register[26][7] ), .D(\register[27][7] ), .S0(n906), .S1(n863), .Y(
        n620) );
  MXI4X1 U1118 ( .A(\register[8][8] ), .B(\register[9][8] ), .C(
        \register[10][8] ), .D(\register[11][8] ), .S0(n908), .S1(n864), .Y(
        n632) );
  MXI4X1 U1119 ( .A(\register[24][8] ), .B(\register[25][8] ), .C(
        \register[26][8] ), .D(\register[27][8] ), .S0(n908), .S1(n864), .Y(
        n628) );
  MXI2X1 U1120 ( .A(n516), .B(n517), .S0(n820), .Y(ReadData2_o[9]) );
  MX4X1 U1121 ( .A(n638), .B(n636), .C(n637), .D(n635), .S0(n826), .S1(n834), 
        .Y(n517) );
  MX4X1 U1122 ( .A(n642), .B(n640), .C(n641), .D(n639), .S0(n826), .S1(n834), 
        .Y(n516) );
  MXI4X1 U1123 ( .A(\register[28][9] ), .B(\register[29][9] ), .C(
        \register[30][9] ), .D(\register[31][9] ), .S0(n908), .S1(n864), .Y(
        n635) );
  MXI2X1 U1124 ( .A(n518), .B(n519), .S0(n820), .Y(ReadData2_o[10]) );
  MX4X1 U1125 ( .A(n646), .B(n644), .C(n645), .D(n643), .S0(n826), .S1(n834), 
        .Y(n519) );
  MX4X1 U1126 ( .A(n650), .B(n648), .C(n649), .D(n647), .S0(n826), .S1(n834), 
        .Y(n518) );
  MXI4X1 U1127 ( .A(\register[28][10] ), .B(\register[29][10] ), .C(
        \register[30][10] ), .D(\register[31][10] ), .S0(n909), .S1(n865), .Y(
        n643) );
  MXI2X1 U1128 ( .A(n520), .B(n521), .S0(n820), .Y(ReadData2_o[11]) );
  MX4X1 U1129 ( .A(n654), .B(n652), .C(n653), .D(n651), .S0(n826), .S1(n834), 
        .Y(n521) );
  MX4X1 U1130 ( .A(n658), .B(n656), .C(n657), .D(n655), .S0(n826), .S1(n834), 
        .Y(n520) );
  MXI4X1 U1131 ( .A(\register[28][11] ), .B(\register[29][11] ), .C(
        \register[30][11] ), .D(\register[31][11] ), .S0(n910), .S1(n866), .Y(
        n651) );
  MXI2X1 U1132 ( .A(n522), .B(n523), .S0(n820), .Y(ReadData2_o[12]) );
  MX4X1 U1133 ( .A(n662), .B(n660), .C(n661), .D(n659), .S0(n826), .S1(n834), 
        .Y(n523) );
  MX4X1 U1134 ( .A(n666), .B(n664), .C(n665), .D(n663), .S0(n826), .S1(n835), 
        .Y(n522) );
  MXI4X1 U1135 ( .A(\register[28][12] ), .B(\register[29][12] ), .C(
        \register[30][12] ), .D(\register[31][12] ), .S0(n910), .S1(n866), .Y(
        n659) );
  MXI2X1 U1136 ( .A(n524), .B(n525), .S0(n820), .Y(ReadData2_o[13]) );
  MX4X1 U1137 ( .A(n670), .B(n668), .C(n669), .D(n667), .S0(n826), .S1(n835), 
        .Y(n525) );
  MX4X1 U1138 ( .A(n674), .B(n672), .C(n673), .D(n671), .S0(n826), .S1(n835), 
        .Y(n524) );
  MXI4X1 U1139 ( .A(\register[28][13] ), .B(\register[29][13] ), .C(
        \register[30][13] ), .D(\register[31][13] ), .S0(n911), .S1(n867), .Y(
        n667) );
  MXI2X1 U1140 ( .A(n526), .B(n527), .S0(n820), .Y(ReadData2_o[14]) );
  MX4X1 U1141 ( .A(n678), .B(n676), .C(n677), .D(n675), .S0(n827), .S1(n835), 
        .Y(n527) );
  MX4X1 U1142 ( .A(n682), .B(n680), .C(n681), .D(n679), .S0(n827), .S1(n835), 
        .Y(n526) );
  MXI4X1 U1143 ( .A(\register[28][14] ), .B(\register[29][14] ), .C(
        \register[30][14] ), .D(\register[31][14] ), .S0(n912), .S1(n868), .Y(
        n675) );
  MXI2X1 U1144 ( .A(n528), .B(n529), .S0(n820), .Y(ReadData2_o[15]) );
  MX4X1 U1145 ( .A(n686), .B(n684), .C(n685), .D(n683), .S0(n827), .S1(n835), 
        .Y(n529) );
  MX4X1 U1146 ( .A(n690), .B(n688), .C(n689), .D(n687), .S0(n827), .S1(n835), 
        .Y(n528) );
  MXI4X1 U1147 ( .A(\register[28][15] ), .B(\register[29][15] ), .C(
        \register[30][15] ), .D(\register[31][15] ), .S0(n912), .S1(n868), .Y(
        n683) );
  MXI2X1 U1148 ( .A(n530), .B(n531), .S0(n820), .Y(ReadData2_o[16]) );
  MX4X1 U1149 ( .A(n694), .B(n692), .C(n693), .D(n691), .S0(n827), .S1(n835), 
        .Y(n531) );
  MX4X1 U1150 ( .A(n698), .B(n696), .C(n697), .D(n695), .S0(n827), .S1(n835), 
        .Y(n530) );
  MXI4X1 U1151 ( .A(\register[28][16] ), .B(\register[29][16] ), .C(
        \register[30][16] ), .D(\register[31][16] ), .S0(n913), .S1(n869), .Y(
        n691) );
  MXI2X1 U1152 ( .A(n532), .B(n533), .S0(n820), .Y(ReadData2_o[17]) );
  MX4X1 U1153 ( .A(n702), .B(n700), .C(n701), .D(n699), .S0(n827), .S1(n835), 
        .Y(n533) );
  MX4X1 U1154 ( .A(n706), .B(n704), .C(n705), .D(n703), .S0(n827), .S1(n835), 
        .Y(n532) );
  MXI4X1 U1155 ( .A(\register[28][17] ), .B(\register[29][17] ), .C(
        \register[30][17] ), .D(\register[31][17] ), .S0(n914), .S1(n870), .Y(
        n699) );
  MXI2X1 U1156 ( .A(n534), .B(n535), .S0(n820), .Y(ReadData2_o[18]) );
  MX4X1 U1157 ( .A(n710), .B(n708), .C(n709), .D(n707), .S0(n827), .S1(n835), 
        .Y(n535) );
  MX4X1 U1158 ( .A(n714), .B(n712), .C(n713), .D(n711), .S0(n827), .S1(n835), 
        .Y(n534) );
  MXI4X1 U1159 ( .A(\register[28][18] ), .B(\register[29][18] ), .C(
        \register[30][18] ), .D(\register[31][18] ), .S0(n914), .S1(n870), .Y(
        n707) );
  MXI2X1 U1160 ( .A(n536), .B(n537), .S0(n820), .Y(ReadData2_o[19]) );
  MX4X1 U1161 ( .A(n718), .B(n716), .C(n717), .D(n715), .S0(n827), .S1(n836), 
        .Y(n537) );
  MX4X1 U1162 ( .A(n722), .B(n720), .C(n721), .D(n719), .S0(n827), .S1(n836), 
        .Y(n536) );
  MXI4X1 U1163 ( .A(\register[28][19] ), .B(\register[29][19] ), .C(
        \register[30][19] ), .D(\register[31][19] ), .S0(n915), .S1(n871), .Y(
        n715) );
  MXI2X1 U1164 ( .A(n538), .B(n539), .S0(n821), .Y(ReadData2_o[20]) );
  MX4X1 U1165 ( .A(n726), .B(n724), .C(n725), .D(n723), .S0(n828), .S1(n836), 
        .Y(n539) );
  MX4X1 U1166 ( .A(n730), .B(n728), .C(n729), .D(n727), .S0(n828), .S1(n836), 
        .Y(n538) );
  MXI4X1 U1167 ( .A(\register[28][20] ), .B(\register[29][20] ), .C(
        \register[30][20] ), .D(\register[31][20] ), .S0(n916), .S1(n874), .Y(
        n723) );
  MXI2X1 U1168 ( .A(n540), .B(n541), .S0(n821), .Y(ReadData2_o[21]) );
  MX4X1 U1169 ( .A(n734), .B(n732), .C(n733), .D(n731), .S0(n828), .S1(n836), 
        .Y(n541) );
  MX4X1 U1170 ( .A(n738), .B(n736), .C(n737), .D(n735), .S0(n828), .S1(n836), 
        .Y(n540) );
  MXI4X1 U1171 ( .A(\register[28][21] ), .B(\register[29][21] ), .C(
        \register[30][21] ), .D(\register[31][21] ), .S0(n916), .S1(n874), .Y(
        n731) );
  MXI2X1 U1172 ( .A(n542), .B(n543), .S0(n821), .Y(ReadData2_o[22]) );
  MX4X1 U1173 ( .A(n742), .B(n740), .C(n741), .D(n739), .S0(n828), .S1(n836), 
        .Y(n543) );
  MX4X1 U1174 ( .A(n746), .B(n744), .C(n745), .D(n743), .S0(n828), .S1(n836), 
        .Y(n542) );
  MXI4X1 U1175 ( .A(\register[28][22] ), .B(\register[29][22] ), .C(
        \register[30][22] ), .D(\register[31][22] ), .S0(n917), .S1(n875), .Y(
        n739) );
  MXI2X1 U1176 ( .A(n544), .B(n545), .S0(n821), .Y(ReadData2_o[23]) );
  MX4X1 U1177 ( .A(n750), .B(n748), .C(n749), .D(n747), .S0(n828), .S1(n836), 
        .Y(n545) );
  MX4X1 U1178 ( .A(n754), .B(n752), .C(n753), .D(n751), .S0(n828), .S1(n836), 
        .Y(n544) );
  MXI4X1 U1179 ( .A(\register[28][23] ), .B(\register[29][23] ), .C(
        \register[30][23] ), .D(\register[31][23] ), .S0(n918), .S1(n876), .Y(
        n747) );
  MXI2X1 U1180 ( .A(n546), .B(n547), .S0(n821), .Y(ReadData2_o[24]) );
  MX4X1 U1181 ( .A(n758), .B(n756), .C(n757), .D(n755), .S0(n828), .S1(n836), 
        .Y(n547) );
  MX4X1 U1182 ( .A(n762), .B(n760), .C(n761), .D(n759), .S0(n828), .S1(n836), 
        .Y(n546) );
  MXI4X1 U1183 ( .A(\register[28][24] ), .B(\register[29][24] ), .C(
        \register[30][24] ), .D(\register[31][24] ), .S0(n918), .S1(n876), .Y(
        n755) );
  MXI2X1 U1184 ( .A(n548), .B(n549), .S0(n821), .Y(ReadData2_o[25]) );
  MX4X1 U1185 ( .A(n766), .B(n764), .C(n765), .D(n763), .S0(n828), .S1(n836), 
        .Y(n549) );
  MX4X1 U1186 ( .A(n770), .B(n768), .C(n769), .D(n767), .S0(n828), .S1(n837), 
        .Y(n548) );
  MXI4X1 U1187 ( .A(\register[28][25] ), .B(\register[29][25] ), .C(
        \register[30][25] ), .D(\register[31][25] ), .S0(n919), .S1(n877), .Y(
        n763) );
  MXI2X1 U1188 ( .A(n550), .B(n551), .S0(n821), .Y(ReadData2_o[26]) );
  MX4X1 U1189 ( .A(n774), .B(n772), .C(n773), .D(n771), .S0(n829), .S1(n837), 
        .Y(n551) );
  MX4X1 U1190 ( .A(n778), .B(n776), .C(n777), .D(n775), .S0(n829), .S1(n837), 
        .Y(n550) );
  MXI4X1 U1191 ( .A(\register[28][26] ), .B(\register[29][26] ), .C(
        \register[30][26] ), .D(\register[31][26] ), .S0(n920), .S1(n878), .Y(
        n771) );
  MXI2X1 U1192 ( .A(n552), .B(n553), .S0(n821), .Y(ReadData2_o[27]) );
  MX4X1 U1193 ( .A(n782), .B(n780), .C(n781), .D(n779), .S0(n829), .S1(n837), 
        .Y(n553) );
  MX4X1 U1194 ( .A(n786), .B(n784), .C(n785), .D(n783), .S0(n829), .S1(n837), 
        .Y(n552) );
  MXI4X1 U1195 ( .A(\register[28][27] ), .B(\register[29][27] ), .C(
        \register[30][27] ), .D(\register[31][27] ), .S0(n920), .S1(n878), .Y(
        n779) );
  MXI2X1 U1196 ( .A(n554), .B(n555), .S0(n821), .Y(ReadData2_o[28]) );
  MX4X1 U1197 ( .A(n790), .B(n788), .C(n789), .D(n787), .S0(n829), .S1(n837), 
        .Y(n555) );
  MX4X1 U1198 ( .A(n794), .B(n792), .C(n793), .D(n791), .S0(n829), .S1(n837), 
        .Y(n554) );
  MXI4X1 U1199 ( .A(\register[28][28] ), .B(\register[29][28] ), .C(
        \register[30][28] ), .D(\register[31][28] ), .S0(n921), .S1(n879), .Y(
        n787) );
  MXI2X1 U1200 ( .A(n556), .B(n557), .S0(n821), .Y(ReadData2_o[29]) );
  MX4X1 U1201 ( .A(n798), .B(n796), .C(n797), .D(n795), .S0(n829), .S1(n837), 
        .Y(n557) );
  MX4X1 U1202 ( .A(n802), .B(n800), .C(n801), .D(n799), .S0(n829), .S1(n837), 
        .Y(n556) );
  MXI4X1 U1203 ( .A(\register[28][29] ), .B(\register[29][29] ), .C(
        \register[30][29] ), .D(\register[31][29] ), .S0(n922), .S1(n880), .Y(
        n795) );
  MXI2X1 U1204 ( .A(n558), .B(n559), .S0(n821), .Y(ReadData2_o[30]) );
  MX4X1 U1205 ( .A(n806), .B(n804), .C(n805), .D(n803), .S0(n829), .S1(n837), 
        .Y(n559) );
  MX4X1 U1206 ( .A(n810), .B(n808), .C(n809), .D(n807), .S0(n829), .S1(n837), 
        .Y(n558) );
  MXI4X1 U1207 ( .A(\register[28][30] ), .B(\register[29][30] ), .C(
        \register[30][30] ), .D(\register[31][30] ), .S0(n922), .S1(n880), .Y(
        n803) );
  MXI2X1 U1208 ( .A(n560), .B(n561), .S0(n821), .Y(ReadData2_o[31]) );
  MX4X1 U1209 ( .A(n814), .B(n812), .C(n813), .D(n811), .S0(n829), .S1(n837), 
        .Y(n561) );
  MX4X1 U1210 ( .A(n818), .B(n816), .C(n817), .D(n815), .S0(n829), .S1(n837), 
        .Y(n560) );
  MXI4X1 U1211 ( .A(\register[28][31] ), .B(\register[29][31] ), .C(
        \register[30][31] ), .D(\register[31][31] ), .S0(n923), .S1(n881), .Y(
        n811) );
  MXI4X1 U1212 ( .A(\register[4][9] ), .B(\register[5][9] ), .C(
        \register[6][9] ), .D(\register[7][9] ), .S0(n909), .S1(n865), .Y(n641) );
  MXI4X1 U1213 ( .A(\register[20][9] ), .B(\register[21][9] ), .C(
        \register[22][9] ), .D(\register[23][9] ), .S0(n908), .S1(n864), .Y(
        n637) );
  MXI4X1 U1214 ( .A(\register[4][10] ), .B(\register[5][10] ), .C(
        \register[6][10] ), .D(\register[7][10] ), .S0(n909), .S1(n865), .Y(
        n649) );
  MXI4X1 U1215 ( .A(\register[20][10] ), .B(\register[21][10] ), .C(
        \register[22][10] ), .D(\register[23][10] ), .S0(n909), .S1(n865), .Y(
        n645) );
  MXI4X1 U1216 ( .A(\register[4][11] ), .B(\register[5][11] ), .C(
        \register[6][11] ), .D(\register[7][11] ), .S0(n910), .S1(n866), .Y(
        n657) );
  MXI4X1 U1217 ( .A(\register[20][11] ), .B(\register[21][11] ), .C(
        \register[22][11] ), .D(\register[23][11] ), .S0(n910), .S1(n866), .Y(
        n653) );
  MXI4X1 U1218 ( .A(\register[4][12] ), .B(\register[5][12] ), .C(
        \register[6][12] ), .D(\register[7][12] ), .S0(n911), .S1(n867), .Y(
        n665) );
  MXI4X1 U1219 ( .A(\register[20][12] ), .B(\register[21][12] ), .C(
        \register[22][12] ), .D(\register[23][12] ), .S0(n910), .S1(n866), .Y(
        n661) );
  MXI4X1 U1220 ( .A(\register[4][13] ), .B(\register[5][13] ), .C(
        \register[6][13] ), .D(\register[7][13] ), .S0(n911), .S1(n867), .Y(
        n673) );
  MXI4X1 U1221 ( .A(\register[20][13] ), .B(\register[21][13] ), .C(
        \register[22][13] ), .D(\register[23][13] ), .S0(n911), .S1(n867), .Y(
        n669) );
  MXI4X1 U1222 ( .A(\register[4][14] ), .B(\register[5][14] ), .C(
        \register[6][14] ), .D(\register[7][14] ), .S0(n912), .S1(n868), .Y(
        n681) );
  MXI4X1 U1223 ( .A(\register[20][14] ), .B(\register[21][14] ), .C(
        \register[22][14] ), .D(\register[23][14] ), .S0(n912), .S1(n868), .Y(
        n677) );
  MXI4X1 U1224 ( .A(\register[4][15] ), .B(\register[5][15] ), .C(
        \register[6][15] ), .D(\register[7][15] ), .S0(n913), .S1(n869), .Y(
        n689) );
  MXI4X1 U1225 ( .A(\register[20][15] ), .B(\register[21][15] ), .C(
        \register[22][15] ), .D(\register[23][15] ), .S0(n912), .S1(n868), .Y(
        n685) );
  MXI4X1 U1226 ( .A(\register[4][16] ), .B(\register[5][16] ), .C(
        \register[6][16] ), .D(\register[7][16] ), .S0(n913), .S1(n869), .Y(
        n697) );
  MXI4X1 U1227 ( .A(\register[20][16] ), .B(\register[21][16] ), .C(
        \register[22][16] ), .D(\register[23][16] ), .S0(n913), .S1(n869), .Y(
        n693) );
  MXI4X1 U1228 ( .A(\register[4][17] ), .B(\register[5][17] ), .C(
        \register[6][17] ), .D(\register[7][17] ), .S0(n914), .S1(n870), .Y(
        n705) );
  MXI4X1 U1229 ( .A(\register[20][17] ), .B(\register[21][17] ), .C(
        \register[22][17] ), .D(\register[23][17] ), .S0(n914), .S1(n870), .Y(
        n701) );
  MXI4X1 U1230 ( .A(\register[4][18] ), .B(\register[5][18] ), .C(
        \register[6][18] ), .D(\register[7][18] ), .S0(n915), .S1(n871), .Y(
        n713) );
  MXI4X1 U1231 ( .A(\register[20][18] ), .B(\register[21][18] ), .C(
        \register[22][18] ), .D(\register[23][18] ), .S0(n914), .S1(n870), .Y(
        n709) );
  MXI4X1 U1232 ( .A(\register[4][19] ), .B(\register[5][19] ), .C(
        \register[6][19] ), .D(\register[7][19] ), .S0(n915), .S1(n871), .Y(
        n721) );
  MXI4X1 U1233 ( .A(\register[20][19] ), .B(\register[21][19] ), .C(
        \register[22][19] ), .D(\register[23][19] ), .S0(n915), .S1(n871), .Y(
        n717) );
  MXI4X1 U1234 ( .A(\register[4][20] ), .B(\register[5][20] ), .C(
        \register[6][20] ), .D(\register[7][20] ), .S0(n916), .S1(n874), .Y(
        n729) );
  MXI4X1 U1235 ( .A(\register[20][20] ), .B(\register[21][20] ), .C(
        \register[22][20] ), .D(\register[23][20] ), .S0(n916), .S1(n874), .Y(
        n725) );
  MXI4X1 U1236 ( .A(\register[4][21] ), .B(\register[5][21] ), .C(
        \register[6][21] ), .D(\register[7][21] ), .S0(n917), .S1(n875), .Y(
        n737) );
  MXI4X1 U1237 ( .A(\register[20][21] ), .B(\register[21][21] ), .C(
        \register[22][21] ), .D(\register[23][21] ), .S0(n916), .S1(n874), .Y(
        n733) );
  MXI4X1 U1238 ( .A(\register[4][22] ), .B(\register[5][22] ), .C(
        \register[6][22] ), .D(\register[7][22] ), .S0(n917), .S1(n875), .Y(
        n745) );
  MXI4X1 U1239 ( .A(\register[20][22] ), .B(\register[21][22] ), .C(
        \register[22][22] ), .D(\register[23][22] ), .S0(n917), .S1(n875), .Y(
        n741) );
  MXI4X1 U1240 ( .A(\register[4][23] ), .B(\register[5][23] ), .C(
        \register[6][23] ), .D(\register[7][23] ), .S0(n918), .S1(n876), .Y(
        n753) );
  MXI4X1 U1241 ( .A(\register[20][23] ), .B(\register[21][23] ), .C(
        \register[22][23] ), .D(\register[23][23] ), .S0(n918), .S1(n876), .Y(
        n749) );
  MXI4X1 U1242 ( .A(\register[4][24] ), .B(\register[5][24] ), .C(
        \register[6][24] ), .D(\register[7][24] ), .S0(n919), .S1(n877), .Y(
        n761) );
  MXI4X1 U1243 ( .A(\register[20][24] ), .B(\register[21][24] ), .C(
        \register[22][24] ), .D(\register[23][24] ), .S0(n918), .S1(n876), .Y(
        n757) );
  MXI4X1 U1244 ( .A(\register[4][25] ), .B(\register[5][25] ), .C(
        \register[6][25] ), .D(\register[7][25] ), .S0(n919), .S1(n877), .Y(
        n769) );
  MXI4X1 U1245 ( .A(\register[20][25] ), .B(\register[21][25] ), .C(
        \register[22][25] ), .D(\register[23][25] ), .S0(n919), .S1(n877), .Y(
        n765) );
  MXI4X1 U1246 ( .A(\register[4][26] ), .B(\register[5][26] ), .C(
        \register[6][26] ), .D(\register[7][26] ), .S0(n920), .S1(n878), .Y(
        n777) );
  MXI4X1 U1247 ( .A(\register[20][26] ), .B(\register[21][26] ), .C(
        \register[22][26] ), .D(\register[23][26] ), .S0(n920), .S1(n878), .Y(
        n773) );
  MXI4X1 U1248 ( .A(\register[4][27] ), .B(\register[5][27] ), .C(
        \register[6][27] ), .D(\register[7][27] ), .S0(n921), .S1(n879), .Y(
        n785) );
  MXI4X1 U1249 ( .A(\register[20][27] ), .B(\register[21][27] ), .C(
        \register[22][27] ), .D(\register[23][27] ), .S0(n920), .S1(n878), .Y(
        n781) );
  MXI4X1 U1250 ( .A(\register[4][28] ), .B(\register[5][28] ), .C(
        \register[6][28] ), .D(\register[7][28] ), .S0(n921), .S1(n879), .Y(
        n793) );
  MXI4X1 U1251 ( .A(\register[20][28] ), .B(\register[21][28] ), .C(
        \register[22][28] ), .D(\register[23][28] ), .S0(n921), .S1(n879), .Y(
        n789) );
  MXI4X1 U1252 ( .A(\register[4][29] ), .B(\register[5][29] ), .C(
        \register[6][29] ), .D(\register[7][29] ), .S0(n922), .S1(n880), .Y(
        n801) );
  MXI4X1 U1253 ( .A(\register[20][29] ), .B(\register[21][29] ), .C(
        \register[22][29] ), .D(\register[23][29] ), .S0(n922), .S1(n880), .Y(
        n797) );
  MXI4X1 U1254 ( .A(\register[4][30] ), .B(\register[5][30] ), .C(
        \register[6][30] ), .D(\register[7][30] ), .S0(n923), .S1(n881), .Y(
        n809) );
  MXI4X1 U1255 ( .A(\register[20][30] ), .B(\register[21][30] ), .C(
        \register[22][30] ), .D(\register[23][30] ), .S0(n922), .S1(n880), .Y(
        n805) );
  MXI4X1 U1256 ( .A(\register[4][31] ), .B(\register[5][31] ), .C(
        \register[6][31] ), .D(\register[7][31] ), .S0(n923), .S1(n881), .Y(
        n817) );
  MXI4X1 U1257 ( .A(\register[20][31] ), .B(\register[21][31] ), .C(
        \register[22][31] ), .D(\register[23][31] ), .S0(n923), .S1(n881), .Y(
        n813) );
  MXI4X1 U1258 ( .A(\register[0][9] ), .B(\register[1][9] ), .C(
        \register[2][9] ), .D(\register[3][9] ), .S0(n909), .S1(n865), .Y(n642) );
  MXI4X1 U1259 ( .A(\register[16][9] ), .B(\register[17][9] ), .C(
        \register[18][9] ), .D(\register[19][9] ), .S0(n908), .S1(n864), .Y(
        n638) );
  MXI4X1 U1260 ( .A(\register[0][10] ), .B(\register[1][10] ), .C(
        \register[2][10] ), .D(\register[3][10] ), .S0(n909), .S1(n865), .Y(
        n650) );
  MXI4X1 U1261 ( .A(\register[16][10] ), .B(\register[17][10] ), .C(
        \register[18][10] ), .D(\register[19][10] ), .S0(n909), .S1(n865), .Y(
        n646) );
  MXI4X1 U1262 ( .A(\register[0][11] ), .B(\register[1][11] ), .C(
        \register[2][11] ), .D(\register[3][11] ), .S0(n910), .S1(n866), .Y(
        n658) );
  MXI4X1 U1263 ( .A(\register[16][11] ), .B(\register[17][11] ), .C(
        \register[18][11] ), .D(\register[19][11] ), .S0(n910), .S1(n866), .Y(
        n654) );
  MXI4X1 U1264 ( .A(\register[0][12] ), .B(\register[1][12] ), .C(
        \register[2][12] ), .D(\register[3][12] ), .S0(n911), .S1(n867), .Y(
        n666) );
  MXI4X1 U1265 ( .A(\register[16][12] ), .B(\register[17][12] ), .C(
        \register[18][12] ), .D(\register[19][12] ), .S0(n910), .S1(n866), .Y(
        n662) );
  MXI4X1 U1266 ( .A(\register[0][13] ), .B(\register[1][13] ), .C(
        \register[2][13] ), .D(\register[3][13] ), .S0(n911), .S1(n867), .Y(
        n674) );
  MXI4X1 U1267 ( .A(\register[16][13] ), .B(\register[17][13] ), .C(
        \register[18][13] ), .D(\register[19][13] ), .S0(n911), .S1(n867), .Y(
        n670) );
  MXI4X1 U1268 ( .A(\register[0][14] ), .B(\register[1][14] ), .C(
        \register[2][14] ), .D(\register[3][14] ), .S0(n912), .S1(n868), .Y(
        n682) );
  MXI4X1 U1269 ( .A(\register[16][14] ), .B(\register[17][14] ), .C(
        \register[18][14] ), .D(\register[19][14] ), .S0(n912), .S1(n868), .Y(
        n678) );
  MXI4X1 U1270 ( .A(\register[0][15] ), .B(\register[1][15] ), .C(
        \register[2][15] ), .D(\register[3][15] ), .S0(n913), .S1(n869), .Y(
        n690) );
  MXI4X1 U1271 ( .A(\register[16][15] ), .B(\register[17][15] ), .C(
        \register[18][15] ), .D(\register[19][15] ), .S0(n912), .S1(n868), .Y(
        n686) );
  MXI4X1 U1272 ( .A(\register[0][16] ), .B(\register[1][16] ), .C(
        \register[2][16] ), .D(\register[3][16] ), .S0(n913), .S1(n869), .Y(
        n698) );
  MXI4X1 U1273 ( .A(\register[16][16] ), .B(\register[17][16] ), .C(
        \register[18][16] ), .D(\register[19][16] ), .S0(n913), .S1(n869), .Y(
        n694) );
  MXI4X1 U1274 ( .A(\register[0][17] ), .B(\register[1][17] ), .C(
        \register[2][17] ), .D(\register[3][17] ), .S0(n914), .S1(n870), .Y(
        n706) );
  MXI4X1 U1275 ( .A(\register[16][17] ), .B(\register[17][17] ), .C(
        \register[18][17] ), .D(\register[19][17] ), .S0(n914), .S1(n870), .Y(
        n702) );
  MXI4X1 U1276 ( .A(\register[0][18] ), .B(\register[1][18] ), .C(
        \register[2][18] ), .D(\register[3][18] ), .S0(n915), .S1(n871), .Y(
        n714) );
  MXI4X1 U1277 ( .A(\register[16][18] ), .B(\register[17][18] ), .C(
        \register[18][18] ), .D(\register[19][18] ), .S0(n914), .S1(n870), .Y(
        n710) );
  MXI4X1 U1278 ( .A(\register[0][19] ), .B(\register[1][19] ), .C(
        \register[2][19] ), .D(\register[3][19] ), .S0(n915), .S1(n871), .Y(
        n722) );
  MXI4X1 U1279 ( .A(\register[16][19] ), .B(\register[17][19] ), .C(
        \register[18][19] ), .D(\register[19][19] ), .S0(n915), .S1(n871), .Y(
        n718) );
  MXI4X1 U1280 ( .A(\register[0][20] ), .B(\register[1][20] ), .C(
        \register[2][20] ), .D(\register[3][20] ), .S0(n916), .S1(n874), .Y(
        n730) );
  MXI4X1 U1281 ( .A(\register[16][20] ), .B(\register[17][20] ), .C(
        \register[18][20] ), .D(\register[19][20] ), .S0(n916), .S1(n874), .Y(
        n726) );
  MXI4X1 U1282 ( .A(\register[0][21] ), .B(\register[1][21] ), .C(
        \register[2][21] ), .D(\register[3][21] ), .S0(n917), .S1(n875), .Y(
        n738) );
  MXI4X1 U1283 ( .A(\register[16][21] ), .B(\register[17][21] ), .C(
        \register[18][21] ), .D(\register[19][21] ), .S0(n916), .S1(n874), .Y(
        n734) );
  MXI4X1 U1284 ( .A(\register[0][22] ), .B(\register[1][22] ), .C(
        \register[2][22] ), .D(\register[3][22] ), .S0(n917), .S1(n875), .Y(
        n746) );
  MXI4X1 U1285 ( .A(\register[16][22] ), .B(\register[17][22] ), .C(
        \register[18][22] ), .D(\register[19][22] ), .S0(n917), .S1(n875), .Y(
        n742) );
  MXI4X1 U1286 ( .A(\register[0][23] ), .B(\register[1][23] ), .C(
        \register[2][23] ), .D(\register[3][23] ), .S0(n918), .S1(n876), .Y(
        n754) );
  MXI4X1 U1287 ( .A(\register[16][23] ), .B(\register[17][23] ), .C(
        \register[18][23] ), .D(\register[19][23] ), .S0(n918), .S1(n876), .Y(
        n750) );
  MXI4X1 U1288 ( .A(\register[0][24] ), .B(\register[1][24] ), .C(
        \register[2][24] ), .D(\register[3][24] ), .S0(n919), .S1(n877), .Y(
        n762) );
  MXI4X1 U1289 ( .A(\register[16][24] ), .B(\register[17][24] ), .C(
        \register[18][24] ), .D(\register[19][24] ), .S0(n918), .S1(n876), .Y(
        n758) );
  MXI4X1 U1290 ( .A(\register[0][25] ), .B(\register[1][25] ), .C(
        \register[2][25] ), .D(\register[3][25] ), .S0(n919), .S1(n877), .Y(
        n770) );
  MXI4X1 U1291 ( .A(\register[16][25] ), .B(\register[17][25] ), .C(
        \register[18][25] ), .D(\register[19][25] ), .S0(n919), .S1(n877), .Y(
        n766) );
  MXI4X1 U1292 ( .A(\register[0][26] ), .B(\register[1][26] ), .C(
        \register[2][26] ), .D(\register[3][26] ), .S0(n920), .S1(n878), .Y(
        n778) );
  MXI4X1 U1293 ( .A(\register[16][26] ), .B(\register[17][26] ), .C(
        \register[18][26] ), .D(\register[19][26] ), .S0(n920), .S1(n878), .Y(
        n774) );
  MXI4X1 U1294 ( .A(\register[0][27] ), .B(\register[1][27] ), .C(
        \register[2][27] ), .D(\register[3][27] ), .S0(n921), .S1(n879), .Y(
        n786) );
  MXI4X1 U1295 ( .A(\register[16][27] ), .B(\register[17][27] ), .C(
        \register[18][27] ), .D(\register[19][27] ), .S0(n920), .S1(n878), .Y(
        n782) );
  MXI4X1 U1296 ( .A(\register[0][28] ), .B(\register[1][28] ), .C(
        \register[2][28] ), .D(\register[3][28] ), .S0(n921), .S1(n879), .Y(
        n794) );
  MXI4X1 U1297 ( .A(\register[16][28] ), .B(\register[17][28] ), .C(
        \register[18][28] ), .D(\register[19][28] ), .S0(n921), .S1(n879), .Y(
        n790) );
  MXI4X1 U1298 ( .A(\register[0][29] ), .B(\register[1][29] ), .C(
        \register[2][29] ), .D(\register[3][29] ), .S0(n922), .S1(n880), .Y(
        n802) );
  MXI4X1 U1299 ( .A(\register[16][29] ), .B(\register[17][29] ), .C(
        \register[18][29] ), .D(\register[19][29] ), .S0(n922), .S1(n880), .Y(
        n798) );
  MXI4X1 U1300 ( .A(\register[0][30] ), .B(\register[1][30] ), .C(
        \register[2][30] ), .D(\register[3][30] ), .S0(n923), .S1(n881), .Y(
        n810) );
  MXI4X1 U1301 ( .A(\register[16][30] ), .B(\register[17][30] ), .C(
        \register[18][30] ), .D(\register[19][30] ), .S0(n922), .S1(n880), .Y(
        n806) );
  MXI4X1 U1302 ( .A(\register[0][31] ), .B(\register[1][31] ), .C(
        \register[2][31] ), .D(\register[3][31] ), .S0(n923), .S1(n881), .Y(
        n818) );
  MXI4X1 U1303 ( .A(\register[16][31] ), .B(\register[17][31] ), .C(
        \register[18][31] ), .D(\register[19][31] ), .S0(n923), .S1(n881), .Y(
        n814) );
  MXI4X1 U1304 ( .A(\register[12][9] ), .B(\register[13][9] ), .C(
        \register[14][9] ), .D(\register[15][9] ), .S0(n909), .S1(n865), .Y(
        n639) );
  MXI4X1 U1305 ( .A(\register[12][10] ), .B(\register[13][10] ), .C(
        \register[14][10] ), .D(\register[15][10] ), .S0(n909), .S1(n865), .Y(
        n647) );
  MXI4X1 U1306 ( .A(\register[12][11] ), .B(\register[13][11] ), .C(
        \register[14][11] ), .D(\register[15][11] ), .S0(n910), .S1(n866), .Y(
        n655) );
  MXI4X1 U1307 ( .A(\register[12][12] ), .B(\register[13][12] ), .C(
        \register[14][12] ), .D(\register[15][12] ), .S0(n911), .S1(n867), .Y(
        n663) );
  MXI4X1 U1308 ( .A(\register[12][13] ), .B(\register[13][13] ), .C(
        \register[14][13] ), .D(\register[15][13] ), .S0(n911), .S1(n867), .Y(
        n671) );
  MXI4X1 U1309 ( .A(\register[12][14] ), .B(\register[13][14] ), .C(
        \register[14][14] ), .D(\register[15][14] ), .S0(n912), .S1(n868), .Y(
        n679) );
  MXI4X1 U1310 ( .A(\register[12][15] ), .B(\register[13][15] ), .C(
        \register[14][15] ), .D(\register[15][15] ), .S0(n913), .S1(n869), .Y(
        n687) );
  MXI4X1 U1311 ( .A(\register[12][16] ), .B(\register[13][16] ), .C(
        \register[14][16] ), .D(\register[15][16] ), .S0(n913), .S1(n869), .Y(
        n695) );
  MXI4X1 U1312 ( .A(\register[12][17] ), .B(\register[13][17] ), .C(
        \register[14][17] ), .D(\register[15][17] ), .S0(n914), .S1(n870), .Y(
        n703) );
  MXI4X1 U1313 ( .A(\register[12][18] ), .B(\register[13][18] ), .C(
        \register[14][18] ), .D(\register[15][18] ), .S0(n915), .S1(n871), .Y(
        n711) );
  MXI4X1 U1314 ( .A(\register[12][19] ), .B(\register[13][19] ), .C(
        \register[14][19] ), .D(\register[15][19] ), .S0(n915), .S1(n871), .Y(
        n719) );
  MXI4X1 U1315 ( .A(\register[12][20] ), .B(\register[13][20] ), .C(
        \register[14][20] ), .D(\register[15][20] ), .S0(n916), .S1(n874), .Y(
        n727) );
  MXI4X1 U1316 ( .A(\register[12][21] ), .B(\register[13][21] ), .C(
        \register[14][21] ), .D(\register[15][21] ), .S0(n917), .S1(n875), .Y(
        n735) );
  MXI4X1 U1317 ( .A(\register[12][22] ), .B(\register[13][22] ), .C(
        \register[14][22] ), .D(\register[15][22] ), .S0(n917), .S1(n875), .Y(
        n743) );
  MXI4X1 U1318 ( .A(\register[12][23] ), .B(\register[13][23] ), .C(
        \register[14][23] ), .D(\register[15][23] ), .S0(n918), .S1(n876), .Y(
        n751) );
  MXI4X1 U1319 ( .A(\register[12][24] ), .B(\register[13][24] ), .C(
        \register[14][24] ), .D(\register[15][24] ), .S0(n919), .S1(n877), .Y(
        n759) );
  MXI4X1 U1320 ( .A(\register[12][25] ), .B(\register[13][25] ), .C(
        \register[14][25] ), .D(\register[15][25] ), .S0(n919), .S1(n877), .Y(
        n767) );
  MXI4X1 U1321 ( .A(\register[12][26] ), .B(\register[13][26] ), .C(
        \register[14][26] ), .D(\register[15][26] ), .S0(n920), .S1(n878), .Y(
        n775) );
  MXI4X1 U1322 ( .A(\register[12][27] ), .B(\register[13][27] ), .C(
        \register[14][27] ), .D(\register[15][27] ), .S0(n921), .S1(n879), .Y(
        n783) );
  MXI4X1 U1323 ( .A(\register[12][28] ), .B(\register[13][28] ), .C(
        \register[14][28] ), .D(\register[15][28] ), .S0(n921), .S1(n879), .Y(
        n791) );
  MXI4X1 U1324 ( .A(\register[12][29] ), .B(\register[13][29] ), .C(
        \register[14][29] ), .D(\register[15][29] ), .S0(n922), .S1(n880), .Y(
        n799) );
  MXI4X1 U1325 ( .A(\register[12][30] ), .B(\register[13][30] ), .C(
        \register[14][30] ), .D(\register[15][30] ), .S0(n923), .S1(n881), .Y(
        n807) );
  MXI4X1 U1326 ( .A(\register[12][31] ), .B(\register[13][31] ), .C(
        \register[14][31] ), .D(\register[15][31] ), .S0(n923), .S1(n881), .Y(
        n815) );
  MXI4X1 U1327 ( .A(\register[8][9] ), .B(\register[9][9] ), .C(
        \register[10][9] ), .D(\register[11][9] ), .S0(n909), .S1(n865), .Y(
        n640) );
  MXI4X1 U1328 ( .A(\register[24][9] ), .B(\register[25][9] ), .C(
        \register[26][9] ), .D(\register[27][9] ), .S0(n908), .S1(n864), .Y(
        n636) );
  MXI4X1 U1329 ( .A(\register[8][10] ), .B(\register[9][10] ), .C(
        \register[10][10] ), .D(\register[11][10] ), .S0(n909), .S1(n865), .Y(
        n648) );
  MXI4X1 U1330 ( .A(\register[24][10] ), .B(\register[25][10] ), .C(
        \register[26][10] ), .D(\register[27][10] ), .S0(n909), .S1(n865), .Y(
        n644) );
  MXI4X1 U1331 ( .A(\register[8][11] ), .B(\register[9][11] ), .C(
        \register[10][11] ), .D(\register[11][11] ), .S0(n910), .S1(n866), .Y(
        n656) );
  MXI4X1 U1332 ( .A(\register[24][11] ), .B(\register[25][11] ), .C(
        \register[26][11] ), .D(\register[27][11] ), .S0(n910), .S1(n866), .Y(
        n652) );
  MXI4X1 U1333 ( .A(\register[8][12] ), .B(\register[9][12] ), .C(
        \register[10][12] ), .D(\register[11][12] ), .S0(n911), .S1(n867), .Y(
        n664) );
  MXI4X1 U1334 ( .A(\register[24][12] ), .B(\register[25][12] ), .C(
        \register[26][12] ), .D(\register[27][12] ), .S0(n910), .S1(n866), .Y(
        n660) );
  MXI4X1 U1335 ( .A(\register[8][13] ), .B(\register[9][13] ), .C(
        \register[10][13] ), .D(\register[11][13] ), .S0(n911), .S1(n867), .Y(
        n672) );
  MXI4X1 U1336 ( .A(\register[24][13] ), .B(\register[25][13] ), .C(
        \register[26][13] ), .D(\register[27][13] ), .S0(n911), .S1(n867), .Y(
        n668) );
  MXI4X1 U1337 ( .A(\register[8][14] ), .B(\register[9][14] ), .C(
        \register[10][14] ), .D(\register[11][14] ), .S0(n912), .S1(n868), .Y(
        n680) );
  MXI4X1 U1338 ( .A(\register[24][14] ), .B(\register[25][14] ), .C(
        \register[26][14] ), .D(\register[27][14] ), .S0(n912), .S1(n868), .Y(
        n676) );
  MXI4X1 U1339 ( .A(\register[8][15] ), .B(\register[9][15] ), .C(
        \register[10][15] ), .D(\register[11][15] ), .S0(n913), .S1(n869), .Y(
        n688) );
  MXI4X1 U1340 ( .A(\register[24][15] ), .B(\register[25][15] ), .C(
        \register[26][15] ), .D(\register[27][15] ), .S0(n912), .S1(n868), .Y(
        n684) );
  MXI4X1 U1341 ( .A(\register[8][16] ), .B(\register[9][16] ), .C(
        \register[10][16] ), .D(\register[11][16] ), .S0(n913), .S1(n869), .Y(
        n696) );
  MXI4X1 U1342 ( .A(\register[24][16] ), .B(\register[25][16] ), .C(
        \register[26][16] ), .D(\register[27][16] ), .S0(n913), .S1(n869), .Y(
        n692) );
  MXI4X1 U1343 ( .A(\register[8][17] ), .B(\register[9][17] ), .C(
        \register[10][17] ), .D(\register[11][17] ), .S0(n914), .S1(n870), .Y(
        n704) );
  MXI4X1 U1344 ( .A(\register[24][17] ), .B(\register[25][17] ), .C(
        \register[26][17] ), .D(\register[27][17] ), .S0(n914), .S1(n870), .Y(
        n700) );
  MXI4X1 U1345 ( .A(\register[8][18] ), .B(\register[9][18] ), .C(
        \register[10][18] ), .D(\register[11][18] ), .S0(n915), .S1(n871), .Y(
        n712) );
  MXI4X1 U1346 ( .A(\register[24][18] ), .B(\register[25][18] ), .C(
        \register[26][18] ), .D(\register[27][18] ), .S0(n914), .S1(n870), .Y(
        n708) );
  MXI4X1 U1347 ( .A(\register[8][19] ), .B(\register[9][19] ), .C(
        \register[10][19] ), .D(\register[11][19] ), .S0(n915), .S1(n871), .Y(
        n720) );
  MXI4X1 U1348 ( .A(\register[24][19] ), .B(\register[25][19] ), .C(
        \register[26][19] ), .D(\register[27][19] ), .S0(n915), .S1(n871), .Y(
        n716) );
  MXI4X1 U1349 ( .A(\register[8][20] ), .B(\register[9][20] ), .C(
        \register[10][20] ), .D(\register[11][20] ), .S0(n916), .S1(n874), .Y(
        n728) );
  MXI4X1 U1350 ( .A(\register[24][20] ), .B(\register[25][20] ), .C(
        \register[26][20] ), .D(\register[27][20] ), .S0(n916), .S1(n874), .Y(
        n724) );
  MXI4X1 U1351 ( .A(\register[8][21] ), .B(\register[9][21] ), .C(
        \register[10][21] ), .D(\register[11][21] ), .S0(n917), .S1(n875), .Y(
        n736) );
  MXI4X1 U1352 ( .A(\register[24][21] ), .B(\register[25][21] ), .C(
        \register[26][21] ), .D(\register[27][21] ), .S0(n916), .S1(n874), .Y(
        n732) );
  MXI4X1 U1353 ( .A(\register[8][22] ), .B(\register[9][22] ), .C(
        \register[10][22] ), .D(\register[11][22] ), .S0(n917), .S1(n875), .Y(
        n744) );
  MXI4X1 U1354 ( .A(\register[24][22] ), .B(\register[25][22] ), .C(
        \register[26][22] ), .D(\register[27][22] ), .S0(n917), .S1(n875), .Y(
        n740) );
  MXI4X1 U1355 ( .A(\register[8][23] ), .B(\register[9][23] ), .C(
        \register[10][23] ), .D(\register[11][23] ), .S0(n918), .S1(n876), .Y(
        n752) );
  MXI4X1 U1356 ( .A(\register[24][23] ), .B(\register[25][23] ), .C(
        \register[26][23] ), .D(\register[27][23] ), .S0(n918), .S1(n876), .Y(
        n748) );
  MXI4X1 U1357 ( .A(\register[8][24] ), .B(\register[9][24] ), .C(
        \register[10][24] ), .D(\register[11][24] ), .S0(n919), .S1(n877), .Y(
        n760) );
  MXI4X1 U1358 ( .A(\register[24][24] ), .B(\register[25][24] ), .C(
        \register[26][24] ), .D(\register[27][24] ), .S0(n918), .S1(n876), .Y(
        n756) );
  MXI4X1 U1359 ( .A(\register[8][25] ), .B(\register[9][25] ), .C(
        \register[10][25] ), .D(\register[11][25] ), .S0(n919), .S1(n877), .Y(
        n768) );
  MXI4X1 U1360 ( .A(\register[24][25] ), .B(\register[25][25] ), .C(
        \register[26][25] ), .D(\register[27][25] ), .S0(n919), .S1(n877), .Y(
        n764) );
  MXI4X1 U1361 ( .A(\register[8][26] ), .B(\register[9][26] ), .C(
        \register[10][26] ), .D(\register[11][26] ), .S0(n920), .S1(n878), .Y(
        n776) );
  MXI4X1 U1362 ( .A(\register[24][26] ), .B(\register[25][26] ), .C(
        \register[26][26] ), .D(\register[27][26] ), .S0(n920), .S1(n878), .Y(
        n772) );
  MXI4X1 U1363 ( .A(\register[8][27] ), .B(\register[9][27] ), .C(
        \register[10][27] ), .D(\register[11][27] ), .S0(n921), .S1(n879), .Y(
        n784) );
  MXI4X1 U1364 ( .A(\register[24][27] ), .B(\register[25][27] ), .C(
        \register[26][27] ), .D(\register[27][27] ), .S0(n920), .S1(n878), .Y(
        n780) );
  MXI4X1 U1365 ( .A(\register[8][28] ), .B(\register[9][28] ), .C(
        \register[10][28] ), .D(\register[11][28] ), .S0(n921), .S1(n879), .Y(
        n792) );
  MXI4X1 U1366 ( .A(\register[24][28] ), .B(\register[25][28] ), .C(
        \register[26][28] ), .D(\register[27][28] ), .S0(n921), .S1(n879), .Y(
        n788) );
  MXI4X1 U1367 ( .A(\register[8][29] ), .B(\register[9][29] ), .C(
        \register[10][29] ), .D(\register[11][29] ), .S0(n922), .S1(n880), .Y(
        n800) );
  MXI4X1 U1368 ( .A(\register[24][29] ), .B(\register[25][29] ), .C(
        \register[26][29] ), .D(\register[27][29] ), .S0(n922), .S1(n880), .Y(
        n796) );
  MXI4X1 U1369 ( .A(\register[8][30] ), .B(\register[9][30] ), .C(
        \register[10][30] ), .D(\register[11][30] ), .S0(n923), .S1(n881), .Y(
        n808) );
  MXI4X1 U1370 ( .A(\register[24][30] ), .B(\register[25][30] ), .C(
        \register[26][30] ), .D(\register[27][30] ), .S0(n922), .S1(n880), .Y(
        n804) );
  MXI4X1 U1371 ( .A(\register[8][31] ), .B(\register[9][31] ), .C(
        \register[10][31] ), .D(\register[11][31] ), .S0(n923), .S1(n881), .Y(
        n816) );
  MXI4X1 U1372 ( .A(\register[24][31] ), .B(\register[25][31] ), .C(
        \register[26][31] ), .D(\register[27][31] ), .S0(n923), .S1(n881), .Y(
        n812) );
  CLKMX2X2 U1373 ( .A(\register[31][7] ), .B(n2085), .S0(n1025), .Y(n2060) );
  CLKMX2X2 U1374 ( .A(\register[30][7] ), .B(n2085), .S0(n1020), .Y(n2028) );
  CLKMX2X2 U1375 ( .A(\register[29][0] ), .B(n1026), .S0(n1017), .Y(n2003) );
  CLKMX2X2 U1376 ( .A(\register[29][7] ), .B(n2085), .S0(n1017), .Y(n1996) );
  CLKMX2X2 U1377 ( .A(\register[28][0] ), .B(n1026), .S0(n1014), .Y(n1971) );
  CLKMX2X2 U1378 ( .A(\register[28][7] ), .B(n2085), .S0(n1014), .Y(n1964) );
  CLKMX2X2 U1379 ( .A(\register[27][7] ), .B(n2085), .S0(n1011), .Y(n1932) );
  CLKMX2X2 U1380 ( .A(\register[26][7] ), .B(n2085), .S0(n1008), .Y(n1900) );
  CLKMX2X2 U1381 ( .A(\register[25][7] ), .B(n2085), .S0(n1005), .Y(n1868) );
  CLKMX2X2 U1382 ( .A(\register[24][7] ), .B(n2085), .S0(n1002), .Y(n1836) );
  CLKMX2X2 U1383 ( .A(\register[23][7] ), .B(n2085), .S0(n999), .Y(n1804) );
  CLKMX2X2 U1384 ( .A(\register[22][7] ), .B(n2085), .S0(n996), .Y(n1772) );
  CLKMX2X2 U1385 ( .A(\register[21][7] ), .B(n2085), .S0(n993), .Y(n1740) );
  CLKMX2X2 U1386 ( .A(\register[20][0] ), .B(n1026), .S0(n990), .Y(n1715) );
  CLKMX2X2 U1387 ( .A(\register[20][7] ), .B(n2085), .S0(n990), .Y(n1708) );
  CLKMX2X2 U1388 ( .A(\register[19][7] ), .B(n2086), .S0(n987), .Y(n1676) );
  CLKMX2X2 U1389 ( .A(\register[18][7] ), .B(n2086), .S0(n984), .Y(n1644) );
  CLKMX2X2 U1390 ( .A(\register[17][7] ), .B(n2086), .S0(n981), .Y(n1612) );
  CLKMX2X2 U1391 ( .A(\register[16][7] ), .B(n2086), .S0(n978), .Y(n1580) );
  CLKMX2X2 U1392 ( .A(\register[15][7] ), .B(n2086), .S0(n974), .Y(n1548) );
  CLKMX2X2 U1393 ( .A(\register[14][7] ), .B(n2086), .S0(n971), .Y(n1516) );
  CLKMX2X2 U1394 ( .A(\register[13][7] ), .B(n2086), .S0(n968), .Y(n1484) );
  CLKMX2X2 U1395 ( .A(\register[12][7] ), .B(n2086), .S0(n965), .Y(n1452) );
  CLKMX2X2 U1396 ( .A(\register[11][7] ), .B(n2086), .S0(n962), .Y(n1420) );
  CLKMX2X2 U1397 ( .A(\register[10][7] ), .B(n2086), .S0(n959), .Y(n1388) );
  CLKMX2X2 U1398 ( .A(\register[9][7] ), .B(n2086), .S0(n956), .Y(n1356) );
  CLKMX2X2 U1399 ( .A(\register[8][7] ), .B(n2086), .S0(n953), .Y(n1324) );
  CLKMX2X2 U1400 ( .A(\register[7][7] ), .B(n2087), .S0(n950), .Y(n1292) );
  CLKMX2X2 U1401 ( .A(\register[6][7] ), .B(n2087), .S0(n947), .Y(n1260) );
  CLKMX2X2 U1402 ( .A(\register[5][7] ), .B(n2087), .S0(n944), .Y(n1228) );
  CLKMX2X2 U1403 ( .A(\register[4][7] ), .B(n2087), .S0(n940), .Y(n1196) );
  CLKMX2X2 U1404 ( .A(\register[3][7] ), .B(n2087), .S0(n937), .Y(n1164) );
  CLKMX2X2 U1405 ( .A(\register[2][7] ), .B(n2087), .S0(n934), .Y(n1132) );
  CLKMX2X2 U1406 ( .A(\register[1][7] ), .B(n2087), .S0(n931), .Y(n1100) );
  CLKMX2X2 U1407 ( .A(\register[0][7] ), .B(n2087), .S0(n928), .Y(n1068) );
  CLKMX2X2 U1408 ( .A(\register[31][8] ), .B(n2090), .S0(n1024), .Y(n2059) );
  CLKMX2X2 U1409 ( .A(\register[31][9] ), .B(n2095), .S0(n1024), .Y(n2058) );
  CLKMX2X2 U1410 ( .A(\register[31][10] ), .B(n2100), .S0(n1024), .Y(n2057) );
  CLKMX2X2 U1411 ( .A(\register[31][11] ), .B(n2105), .S0(n1024), .Y(n2056) );
  CLKMX2X2 U1412 ( .A(\register[31][12] ), .B(n2110), .S0(n1024), .Y(n2055) );
  CLKMX2X2 U1413 ( .A(\register[31][13] ), .B(n2115), .S0(n1024), .Y(n2054) );
  CLKMX2X2 U1414 ( .A(\register[31][14] ), .B(n2120), .S0(n1024), .Y(n2053) );
  CLKMX2X2 U1415 ( .A(\register[31][15] ), .B(n2125), .S0(n1024), .Y(n2052) );
  CLKMX2X2 U1416 ( .A(\register[31][16] ), .B(n2130), .S0(n1024), .Y(n2051) );
  CLKMX2X2 U1417 ( .A(\register[31][17] ), .B(n2135), .S0(n1024), .Y(n2050) );
  CLKMX2X2 U1418 ( .A(\register[31][18] ), .B(n2140), .S0(n1024), .Y(n2049) );
  CLKMX2X2 U1419 ( .A(\register[31][19] ), .B(n2145), .S0(n1024), .Y(n2048) );
  CLKMX2X2 U1420 ( .A(\register[31][20] ), .B(n2150), .S0(n1023), .Y(n2047) );
  CLKMX2X2 U1421 ( .A(\register[31][21] ), .B(n2155), .S0(n1023), .Y(n2046) );
  CLKMX2X2 U1422 ( .A(\register[31][22] ), .B(n2160), .S0(n1023), .Y(n2045) );
  CLKMX2X2 U1423 ( .A(\register[31][23] ), .B(n2165), .S0(n1023), .Y(n2044) );
  CLKMX2X2 U1424 ( .A(\register[31][24] ), .B(n2170), .S0(n1023), .Y(n2043) );
  CLKMX2X2 U1425 ( .A(\register[31][25] ), .B(n2175), .S0(n1023), .Y(n2042) );
  CLKMX2X2 U1426 ( .A(\register[31][26] ), .B(n2180), .S0(n1023), .Y(n2041) );
  CLKMX2X2 U1427 ( .A(\register[31][27] ), .B(n2185), .S0(n1023), .Y(n2040) );
  CLKMX2X2 U1428 ( .A(\register[31][28] ), .B(n2190), .S0(n1023), .Y(n2039) );
  CLKMX2X2 U1429 ( .A(\register[31][29] ), .B(n2195), .S0(n1023), .Y(n2038) );
  CLKMX2X2 U1430 ( .A(\register[31][30] ), .B(n2200), .S0(n1023), .Y(n2037) );
  CLKMX2X2 U1431 ( .A(\register[31][31] ), .B(n2205), .S0(n1023), .Y(n2036) );
  CLKMX2X2 U1432 ( .A(\register[30][8] ), .B(n2090), .S0(n1019), .Y(n2027) );
  CLKMX2X2 U1433 ( .A(\register[30][9] ), .B(n2095), .S0(n1019), .Y(n2026) );
  CLKMX2X2 U1434 ( .A(\register[30][10] ), .B(n2100), .S0(n1019), .Y(n2025) );
  CLKMX2X2 U1435 ( .A(\register[30][11] ), .B(n2105), .S0(n1019), .Y(n2024) );
  CLKMX2X2 U1436 ( .A(\register[30][12] ), .B(n2110), .S0(n1019), .Y(n2023) );
  CLKMX2X2 U1437 ( .A(\register[30][13] ), .B(n2115), .S0(n1019), .Y(n2022) );
  CLKMX2X2 U1438 ( .A(\register[30][14] ), .B(n2120), .S0(n1019), .Y(n2021) );
  CLKMX2X2 U1439 ( .A(\register[30][15] ), .B(n2125), .S0(n1019), .Y(n2020) );
  CLKMX2X2 U1440 ( .A(\register[30][16] ), .B(n2130), .S0(n1019), .Y(n2019) );
  CLKMX2X2 U1441 ( .A(\register[30][17] ), .B(n2135), .S0(n1019), .Y(n2018) );
  CLKMX2X2 U1442 ( .A(\register[30][18] ), .B(n2140), .S0(n1019), .Y(n2017) );
  CLKMX2X2 U1443 ( .A(\register[30][19] ), .B(n2145), .S0(n1019), .Y(n2016) );
  CLKMX2X2 U1444 ( .A(\register[30][20] ), .B(n2150), .S0(n1018), .Y(n2015) );
  CLKMX2X2 U1445 ( .A(\register[30][21] ), .B(n2155), .S0(n1018), .Y(n2014) );
  CLKMX2X2 U1446 ( .A(\register[30][22] ), .B(n2160), .S0(n1018), .Y(n2013) );
  CLKMX2X2 U1447 ( .A(\register[30][23] ), .B(n2165), .S0(n1018), .Y(n2012) );
  CLKMX2X2 U1448 ( .A(\register[30][24] ), .B(n2170), .S0(n1018), .Y(n2011) );
  CLKMX2X2 U1449 ( .A(\register[30][25] ), .B(n2175), .S0(n1018), .Y(n2010) );
  CLKMX2X2 U1450 ( .A(\register[30][26] ), .B(n2180), .S0(n1018), .Y(n2009) );
  CLKMX2X2 U1451 ( .A(\register[30][27] ), .B(n2185), .S0(n1018), .Y(n2008) );
  CLKMX2X2 U1452 ( .A(\register[30][28] ), .B(n2190), .S0(n1018), .Y(n2007) );
  CLKMX2X2 U1453 ( .A(\register[30][29] ), .B(n2195), .S0(n1018), .Y(n2006) );
  CLKMX2X2 U1454 ( .A(\register[30][30] ), .B(n2200), .S0(n1018), .Y(n2005) );
  CLKMX2X2 U1455 ( .A(\register[30][31] ), .B(n2205), .S0(n1018), .Y(n2004) );
  CLKMX2X2 U1456 ( .A(\register[29][8] ), .B(n2090), .S0(n1016), .Y(n1995) );
  CLKMX2X2 U1457 ( .A(\register[29][9] ), .B(n2095), .S0(n1016), .Y(n1994) );
  CLKMX2X2 U1458 ( .A(\register[29][10] ), .B(n2100), .S0(n1016), .Y(n1993) );
  CLKMX2X2 U1459 ( .A(\register[29][11] ), .B(n2105), .S0(n1016), .Y(n1992) );
  CLKMX2X2 U1460 ( .A(\register[29][12] ), .B(n2110), .S0(n1016), .Y(n1991) );
  CLKMX2X2 U1461 ( .A(\register[29][13] ), .B(n2115), .S0(n1016), .Y(n1990) );
  CLKMX2X2 U1462 ( .A(\register[29][14] ), .B(n2120), .S0(n1016), .Y(n1989) );
  CLKMX2X2 U1463 ( .A(\register[29][15] ), .B(n2125), .S0(n1016), .Y(n1988) );
  CLKMX2X2 U1464 ( .A(\register[29][16] ), .B(n2130), .S0(n1016), .Y(n1987) );
  CLKMX2X2 U1465 ( .A(\register[29][17] ), .B(n2135), .S0(n1016), .Y(n1986) );
  CLKMX2X2 U1466 ( .A(\register[29][18] ), .B(n2140), .S0(n1016), .Y(n1985) );
  CLKMX2X2 U1467 ( .A(\register[29][19] ), .B(n2145), .S0(n1016), .Y(n1984) );
  CLKMX2X2 U1468 ( .A(\register[29][20] ), .B(n2150), .S0(n1015), .Y(n1983) );
  CLKMX2X2 U1469 ( .A(\register[29][21] ), .B(n2155), .S0(n1015), .Y(n1982) );
  CLKMX2X2 U1470 ( .A(\register[29][22] ), .B(n2160), .S0(n1015), .Y(n1981) );
  CLKMX2X2 U1471 ( .A(\register[29][23] ), .B(n2165), .S0(n1015), .Y(n1980) );
  CLKMX2X2 U1472 ( .A(\register[29][24] ), .B(n2170), .S0(n1015), .Y(n1979) );
  CLKMX2X2 U1473 ( .A(\register[29][25] ), .B(n2175), .S0(n1015), .Y(n1978) );
  CLKMX2X2 U1474 ( .A(\register[29][26] ), .B(n2180), .S0(n1015), .Y(n1977) );
  CLKMX2X2 U1475 ( .A(\register[29][27] ), .B(n2185), .S0(n1015), .Y(n1976) );
  CLKMX2X2 U1476 ( .A(\register[29][28] ), .B(n2190), .S0(n1015), .Y(n1975) );
  CLKMX2X2 U1477 ( .A(\register[29][29] ), .B(n2195), .S0(n1015), .Y(n1974) );
  CLKMX2X2 U1478 ( .A(\register[29][30] ), .B(n2200), .S0(n1015), .Y(n1973) );
  CLKMX2X2 U1479 ( .A(\register[29][31] ), .B(n2205), .S0(n1015), .Y(n1972) );
  CLKMX2X2 U1480 ( .A(\register[28][8] ), .B(n2090), .S0(n1013), .Y(n1963) );
  CLKMX2X2 U1481 ( .A(\register[28][9] ), .B(n2095), .S0(n1013), .Y(n1962) );
  CLKMX2X2 U1482 ( .A(\register[28][10] ), .B(n2100), .S0(n1013), .Y(n1961) );
  CLKMX2X2 U1483 ( .A(\register[28][11] ), .B(n2105), .S0(n1013), .Y(n1960) );
  CLKMX2X2 U1484 ( .A(\register[28][12] ), .B(n2110), .S0(n1013), .Y(n1959) );
  CLKMX2X2 U1485 ( .A(\register[28][13] ), .B(n2115), .S0(n1013), .Y(n1958) );
  CLKMX2X2 U1486 ( .A(\register[28][14] ), .B(n2120), .S0(n1013), .Y(n1957) );
  CLKMX2X2 U1487 ( .A(\register[28][15] ), .B(n2125), .S0(n1013), .Y(n1956) );
  CLKMX2X2 U1488 ( .A(\register[28][16] ), .B(n2130), .S0(n1013), .Y(n1955) );
  CLKMX2X2 U1489 ( .A(\register[28][17] ), .B(n2135), .S0(n1013), .Y(n1954) );
  CLKMX2X2 U1490 ( .A(\register[28][18] ), .B(n2140), .S0(n1013), .Y(n1953) );
  CLKMX2X2 U1491 ( .A(\register[28][19] ), .B(n2145), .S0(n1013), .Y(n1952) );
  CLKMX2X2 U1492 ( .A(\register[28][20] ), .B(n2150), .S0(n1012), .Y(n1951) );
  CLKMX2X2 U1493 ( .A(\register[28][21] ), .B(n2155), .S0(n1012), .Y(n1950) );
  CLKMX2X2 U1494 ( .A(\register[28][22] ), .B(n2160), .S0(n1012), .Y(n1949) );
  CLKMX2X2 U1495 ( .A(\register[28][23] ), .B(n2165), .S0(n1012), .Y(n1948) );
  CLKMX2X2 U1496 ( .A(\register[28][24] ), .B(n2170), .S0(n1012), .Y(n1947) );
  CLKMX2X2 U1497 ( .A(\register[28][25] ), .B(n2175), .S0(n1012), .Y(n1946) );
  CLKMX2X2 U1498 ( .A(\register[28][26] ), .B(n2180), .S0(n1012), .Y(n1945) );
  CLKMX2X2 U1499 ( .A(\register[28][27] ), .B(n2185), .S0(n1012), .Y(n1944) );
  CLKMX2X2 U1500 ( .A(\register[28][28] ), .B(n2190), .S0(n1012), .Y(n1943) );
  CLKMX2X2 U1501 ( .A(\register[28][29] ), .B(n2195), .S0(n1012), .Y(n1942) );
  CLKMX2X2 U1502 ( .A(\register[28][30] ), .B(n2200), .S0(n1012), .Y(n1941) );
  CLKMX2X2 U1503 ( .A(\register[28][31] ), .B(n2205), .S0(n1012), .Y(n1940) );
  CLKMX2X2 U1504 ( .A(\register[27][8] ), .B(n2090), .S0(n1010), .Y(n1931) );
  CLKMX2X2 U1505 ( .A(\register[27][9] ), .B(n2095), .S0(n1010), .Y(n1930) );
  CLKMX2X2 U1506 ( .A(\register[27][10] ), .B(n2100), .S0(n1010), .Y(n1929) );
  CLKMX2X2 U1507 ( .A(\register[27][11] ), .B(n2105), .S0(n1010), .Y(n1928) );
  CLKMX2X2 U1508 ( .A(\register[27][12] ), .B(n2110), .S0(n1010), .Y(n1927) );
  CLKMX2X2 U1509 ( .A(\register[27][13] ), .B(n2115), .S0(n1010), .Y(n1926) );
  CLKMX2X2 U1510 ( .A(\register[27][14] ), .B(n2120), .S0(n1010), .Y(n1925) );
  CLKMX2X2 U1511 ( .A(\register[27][15] ), .B(n2125), .S0(n1010), .Y(n1924) );
  CLKMX2X2 U1512 ( .A(\register[27][16] ), .B(n2130), .S0(n1010), .Y(n1923) );
  CLKMX2X2 U1513 ( .A(\register[27][17] ), .B(n2135), .S0(n1010), .Y(n1922) );
  CLKMX2X2 U1514 ( .A(\register[27][18] ), .B(n2140), .S0(n1010), .Y(n1921) );
  CLKMX2X2 U1515 ( .A(\register[27][19] ), .B(n2145), .S0(n1010), .Y(n1920) );
  CLKMX2X2 U1516 ( .A(\register[27][20] ), .B(n2150), .S0(n1009), .Y(n1919) );
  CLKMX2X2 U1517 ( .A(\register[27][21] ), .B(n2155), .S0(n1009), .Y(n1918) );
  CLKMX2X2 U1518 ( .A(\register[27][22] ), .B(n2160), .S0(n1009), .Y(n1917) );
  CLKMX2X2 U1519 ( .A(\register[27][23] ), .B(n2165), .S0(n1009), .Y(n1916) );
  CLKMX2X2 U1520 ( .A(\register[27][24] ), .B(n2170), .S0(n1009), .Y(n1915) );
  CLKMX2X2 U1521 ( .A(\register[27][25] ), .B(n2175), .S0(n1009), .Y(n1914) );
  CLKMX2X2 U1522 ( .A(\register[27][26] ), .B(n2180), .S0(n1009), .Y(n1913) );
  CLKMX2X2 U1523 ( .A(\register[27][27] ), .B(n2185), .S0(n1009), .Y(n1912) );
  CLKMX2X2 U1524 ( .A(\register[27][28] ), .B(n2190), .S0(n1009), .Y(n1911) );
  CLKMX2X2 U1525 ( .A(\register[27][29] ), .B(n2195), .S0(n1009), .Y(n1910) );
  CLKMX2X2 U1526 ( .A(\register[27][30] ), .B(n2200), .S0(n1009), .Y(n1909) );
  CLKMX2X2 U1527 ( .A(\register[27][31] ), .B(n2205), .S0(n1009), .Y(n1908) );
  CLKMX2X2 U1528 ( .A(\register[26][8] ), .B(n2090), .S0(n1007), .Y(n1899) );
  CLKMX2X2 U1529 ( .A(\register[26][9] ), .B(n2095), .S0(n1007), .Y(n1898) );
  CLKMX2X2 U1530 ( .A(\register[26][10] ), .B(n2100), .S0(n1007), .Y(n1897) );
  CLKMX2X2 U1531 ( .A(\register[26][11] ), .B(n2105), .S0(n1007), .Y(n1896) );
  CLKMX2X2 U1532 ( .A(\register[26][12] ), .B(n2110), .S0(n1007), .Y(n1895) );
  CLKMX2X2 U1533 ( .A(\register[26][13] ), .B(n2115), .S0(n1007), .Y(n1894) );
  CLKMX2X2 U1534 ( .A(\register[26][14] ), .B(n2120), .S0(n1007), .Y(n1893) );
  CLKMX2X2 U1535 ( .A(\register[26][15] ), .B(n2125), .S0(n1007), .Y(n1892) );
  CLKMX2X2 U1536 ( .A(\register[26][16] ), .B(n2130), .S0(n1007), .Y(n1891) );
  CLKMX2X2 U1537 ( .A(\register[26][17] ), .B(n2135), .S0(n1007), .Y(n1890) );
  CLKMX2X2 U1538 ( .A(\register[26][18] ), .B(n2140), .S0(n1007), .Y(n1889) );
  CLKMX2X2 U1539 ( .A(\register[26][19] ), .B(n2145), .S0(n1007), .Y(n1888) );
  CLKMX2X2 U1540 ( .A(\register[26][20] ), .B(n2150), .S0(n1006), .Y(n1887) );
  CLKMX2X2 U1541 ( .A(\register[26][21] ), .B(n2155), .S0(n1006), .Y(n1886) );
  CLKMX2X2 U1542 ( .A(\register[26][22] ), .B(n2160), .S0(n1006), .Y(n1885) );
  CLKMX2X2 U1543 ( .A(\register[26][23] ), .B(n2165), .S0(n1006), .Y(n1884) );
  CLKMX2X2 U1544 ( .A(\register[26][24] ), .B(n2170), .S0(n1006), .Y(n1883) );
  CLKMX2X2 U1545 ( .A(\register[26][25] ), .B(n2175), .S0(n1006), .Y(n1882) );
  CLKMX2X2 U1546 ( .A(\register[26][26] ), .B(n2180), .S0(n1006), .Y(n1881) );
  CLKMX2X2 U1547 ( .A(\register[26][27] ), .B(n2185), .S0(n1006), .Y(n1880) );
  CLKMX2X2 U1548 ( .A(\register[26][28] ), .B(n2190), .S0(n1006), .Y(n1879) );
  CLKMX2X2 U1549 ( .A(\register[26][29] ), .B(n2195), .S0(n1006), .Y(n1878) );
  CLKMX2X2 U1550 ( .A(\register[26][30] ), .B(n2200), .S0(n1006), .Y(n1877) );
  CLKMX2X2 U1551 ( .A(\register[26][31] ), .B(n2205), .S0(n1006), .Y(n1876) );
  CLKMX2X2 U1552 ( .A(\register[25][8] ), .B(n2090), .S0(n1004), .Y(n1867) );
  CLKMX2X2 U1553 ( .A(\register[25][9] ), .B(n2095), .S0(n1004), .Y(n1866) );
  CLKMX2X2 U1554 ( .A(\register[25][10] ), .B(n2100), .S0(n1004), .Y(n1865) );
  CLKMX2X2 U1555 ( .A(\register[25][11] ), .B(n2105), .S0(n1004), .Y(n1864) );
  CLKMX2X2 U1556 ( .A(\register[25][12] ), .B(n2110), .S0(n1004), .Y(n1863) );
  CLKMX2X2 U1557 ( .A(\register[25][13] ), .B(n2115), .S0(n1004), .Y(n1862) );
  CLKMX2X2 U1558 ( .A(\register[25][14] ), .B(n2120), .S0(n1004), .Y(n1861) );
  CLKMX2X2 U1559 ( .A(\register[25][15] ), .B(n2125), .S0(n1004), .Y(n1860) );
  CLKMX2X2 U1560 ( .A(\register[25][16] ), .B(n2130), .S0(n1004), .Y(n1859) );
  CLKMX2X2 U1561 ( .A(\register[25][17] ), .B(n2135), .S0(n1004), .Y(n1858) );
  CLKMX2X2 U1562 ( .A(\register[25][18] ), .B(n2140), .S0(n1004), .Y(n1857) );
  CLKMX2X2 U1563 ( .A(\register[25][19] ), .B(n2145), .S0(n1004), .Y(n1856) );
  CLKMX2X2 U1564 ( .A(\register[25][20] ), .B(n2150), .S0(n1003), .Y(n1855) );
  CLKMX2X2 U1565 ( .A(\register[25][21] ), .B(n2155), .S0(n1003), .Y(n1854) );
  CLKMX2X2 U1566 ( .A(\register[25][22] ), .B(n2160), .S0(n1003), .Y(n1853) );
  CLKMX2X2 U1567 ( .A(\register[25][23] ), .B(n2165), .S0(n1003), .Y(n1852) );
  CLKMX2X2 U1568 ( .A(\register[25][24] ), .B(n2170), .S0(n1003), .Y(n1851) );
  CLKMX2X2 U1569 ( .A(\register[25][25] ), .B(n2175), .S0(n1003), .Y(n1850) );
  CLKMX2X2 U1570 ( .A(\register[25][26] ), .B(n2180), .S0(n1003), .Y(n1849) );
  CLKMX2X2 U1571 ( .A(\register[25][27] ), .B(n2185), .S0(n1003), .Y(n1848) );
  CLKMX2X2 U1572 ( .A(\register[25][28] ), .B(n2190), .S0(n1003), .Y(n1847) );
  CLKMX2X2 U1573 ( .A(\register[25][29] ), .B(n2195), .S0(n1003), .Y(n1846) );
  CLKMX2X2 U1574 ( .A(\register[25][30] ), .B(n2200), .S0(n1003), .Y(n1845) );
  CLKMX2X2 U1575 ( .A(\register[25][31] ), .B(n2205), .S0(n1003), .Y(n1844) );
  CLKMX2X2 U1576 ( .A(\register[24][8] ), .B(n2090), .S0(n1001), .Y(n1835) );
  CLKMX2X2 U1577 ( .A(\register[24][9] ), .B(n2095), .S0(n1001), .Y(n1834) );
  CLKMX2X2 U1578 ( .A(\register[24][10] ), .B(n2100), .S0(n1001), .Y(n1833) );
  CLKMX2X2 U1579 ( .A(\register[24][11] ), .B(n2105), .S0(n1001), .Y(n1832) );
  CLKMX2X2 U1580 ( .A(\register[24][12] ), .B(n2110), .S0(n1001), .Y(n1831) );
  CLKMX2X2 U1581 ( .A(\register[24][13] ), .B(n2115), .S0(n1001), .Y(n1830) );
  CLKMX2X2 U1582 ( .A(\register[24][14] ), .B(n2120), .S0(n1001), .Y(n1829) );
  CLKMX2X2 U1583 ( .A(\register[24][15] ), .B(n2125), .S0(n1001), .Y(n1828) );
  CLKMX2X2 U1584 ( .A(\register[24][16] ), .B(n2130), .S0(n1001), .Y(n1827) );
  CLKMX2X2 U1585 ( .A(\register[24][17] ), .B(n2135), .S0(n1001), .Y(n1826) );
  CLKMX2X2 U1586 ( .A(\register[24][18] ), .B(n2140), .S0(n1001), .Y(n1825) );
  CLKMX2X2 U1587 ( .A(\register[24][19] ), .B(n2145), .S0(n1001), .Y(n1824) );
  CLKMX2X2 U1588 ( .A(\register[24][20] ), .B(n2150), .S0(n1000), .Y(n1823) );
  CLKMX2X2 U1589 ( .A(\register[24][21] ), .B(n2155), .S0(n1000), .Y(n1822) );
  CLKMX2X2 U1590 ( .A(\register[24][22] ), .B(n2160), .S0(n1000), .Y(n1821) );
  CLKMX2X2 U1591 ( .A(\register[24][23] ), .B(n2165), .S0(n1000), .Y(n1820) );
  CLKMX2X2 U1592 ( .A(\register[24][24] ), .B(n2170), .S0(n1000), .Y(n1819) );
  CLKMX2X2 U1593 ( .A(\register[24][25] ), .B(n2175), .S0(n1000), .Y(n1818) );
  CLKMX2X2 U1594 ( .A(\register[24][26] ), .B(n2180), .S0(n1000), .Y(n1817) );
  CLKMX2X2 U1595 ( .A(\register[24][27] ), .B(n2185), .S0(n1000), .Y(n1816) );
  CLKMX2X2 U1596 ( .A(\register[24][28] ), .B(n2190), .S0(n1000), .Y(n1815) );
  CLKMX2X2 U1597 ( .A(\register[24][29] ), .B(n2195), .S0(n1000), .Y(n1814) );
  CLKMX2X2 U1598 ( .A(\register[24][30] ), .B(n2200), .S0(n1000), .Y(n1813) );
  CLKMX2X2 U1599 ( .A(\register[24][31] ), .B(n2205), .S0(n1000), .Y(n1812) );
  CLKMX2X2 U1600 ( .A(\register[23][8] ), .B(n2090), .S0(n998), .Y(n1803) );
  CLKMX2X2 U1601 ( .A(\register[23][9] ), .B(n2095), .S0(n998), .Y(n1802) );
  CLKMX2X2 U1602 ( .A(\register[23][10] ), .B(n2100), .S0(n998), .Y(n1801) );
  CLKMX2X2 U1603 ( .A(\register[23][11] ), .B(n2105), .S0(n998), .Y(n1800) );
  CLKMX2X2 U1604 ( .A(\register[23][12] ), .B(n2110), .S0(n998), .Y(n1799) );
  CLKMX2X2 U1605 ( .A(\register[23][13] ), .B(n2115), .S0(n998), .Y(n1798) );
  CLKMX2X2 U1606 ( .A(\register[23][14] ), .B(n2120), .S0(n998), .Y(n1797) );
  CLKMX2X2 U1607 ( .A(\register[23][15] ), .B(n2125), .S0(n998), .Y(n1796) );
  CLKMX2X2 U1608 ( .A(\register[23][16] ), .B(n2130), .S0(n998), .Y(n1795) );
  CLKMX2X2 U1609 ( .A(\register[23][17] ), .B(n2135), .S0(n998), .Y(n1794) );
  CLKMX2X2 U1610 ( .A(\register[23][18] ), .B(n2140), .S0(n998), .Y(n1793) );
  CLKMX2X2 U1611 ( .A(\register[23][19] ), .B(n2145), .S0(n998), .Y(n1792) );
  CLKMX2X2 U1612 ( .A(\register[23][20] ), .B(n2150), .S0(n997), .Y(n1791) );
  CLKMX2X2 U1613 ( .A(\register[23][21] ), .B(n2155), .S0(n997), .Y(n1790) );
  CLKMX2X2 U1614 ( .A(\register[23][22] ), .B(n2160), .S0(n997), .Y(n1789) );
  CLKMX2X2 U1615 ( .A(\register[23][23] ), .B(n2165), .S0(n997), .Y(n1788) );
  CLKMX2X2 U1616 ( .A(\register[23][24] ), .B(n2170), .S0(n997), .Y(n1787) );
  CLKMX2X2 U1617 ( .A(\register[23][25] ), .B(n2175), .S0(n997), .Y(n1786) );
  CLKMX2X2 U1618 ( .A(\register[23][26] ), .B(n2180), .S0(n997), .Y(n1785) );
  CLKMX2X2 U1619 ( .A(\register[23][27] ), .B(n2185), .S0(n997), .Y(n1784) );
  CLKMX2X2 U1620 ( .A(\register[23][28] ), .B(n2190), .S0(n997), .Y(n1783) );
  CLKMX2X2 U1621 ( .A(\register[23][29] ), .B(n2195), .S0(n997), .Y(n1782) );
  CLKMX2X2 U1622 ( .A(\register[23][30] ), .B(n2200), .S0(n997), .Y(n1781) );
  CLKMX2X2 U1623 ( .A(\register[23][31] ), .B(n2205), .S0(n997), .Y(n1780) );
  CLKMX2X2 U1624 ( .A(\register[22][8] ), .B(n2090), .S0(n995), .Y(n1771) );
  CLKMX2X2 U1625 ( .A(\register[22][9] ), .B(n2095), .S0(n995), .Y(n1770) );
  CLKMX2X2 U1626 ( .A(\register[22][10] ), .B(n2100), .S0(n995), .Y(n1769) );
  CLKMX2X2 U1627 ( .A(\register[22][11] ), .B(n2105), .S0(n995), .Y(n1768) );
  CLKMX2X2 U1628 ( .A(\register[22][12] ), .B(n2110), .S0(n995), .Y(n1767) );
  CLKMX2X2 U1629 ( .A(\register[22][13] ), .B(n2115), .S0(n995), .Y(n1766) );
  CLKMX2X2 U1630 ( .A(\register[22][14] ), .B(n2120), .S0(n995), .Y(n1765) );
  CLKMX2X2 U1631 ( .A(\register[22][15] ), .B(n2125), .S0(n995), .Y(n1764) );
  CLKMX2X2 U1632 ( .A(\register[22][16] ), .B(n2130), .S0(n995), .Y(n1763) );
  CLKMX2X2 U1633 ( .A(\register[22][17] ), .B(n2135), .S0(n995), .Y(n1762) );
  CLKMX2X2 U1634 ( .A(\register[22][18] ), .B(n2140), .S0(n995), .Y(n1761) );
  CLKMX2X2 U1635 ( .A(\register[22][19] ), .B(n2145), .S0(n995), .Y(n1760) );
  CLKMX2X2 U1636 ( .A(\register[22][20] ), .B(n2150), .S0(n994), .Y(n1759) );
  CLKMX2X2 U1637 ( .A(\register[22][21] ), .B(n2155), .S0(n994), .Y(n1758) );
  CLKMX2X2 U1638 ( .A(\register[22][22] ), .B(n2160), .S0(n994), .Y(n1757) );
  CLKMX2X2 U1639 ( .A(\register[22][23] ), .B(n2165), .S0(n994), .Y(n1756) );
  CLKMX2X2 U1640 ( .A(\register[22][24] ), .B(n2170), .S0(n994), .Y(n1755) );
  CLKMX2X2 U1641 ( .A(\register[22][25] ), .B(n2175), .S0(n994), .Y(n1754) );
  CLKMX2X2 U1642 ( .A(\register[22][26] ), .B(n2180), .S0(n994), .Y(n1753) );
  CLKMX2X2 U1643 ( .A(\register[22][27] ), .B(n2185), .S0(n994), .Y(n1752) );
  CLKMX2X2 U1644 ( .A(\register[22][28] ), .B(n2190), .S0(n994), .Y(n1751) );
  CLKMX2X2 U1645 ( .A(\register[22][29] ), .B(n2195), .S0(n994), .Y(n1750) );
  CLKMX2X2 U1646 ( .A(\register[22][30] ), .B(n2200), .S0(n994), .Y(n1749) );
  CLKMX2X2 U1647 ( .A(\register[22][31] ), .B(n2205), .S0(n994), .Y(n1748) );
  CLKMX2X2 U1648 ( .A(\register[21][8] ), .B(n2090), .S0(n992), .Y(n1739) );
  CLKMX2X2 U1649 ( .A(\register[21][9] ), .B(n2095), .S0(n992), .Y(n1738) );
  CLKMX2X2 U1650 ( .A(\register[21][10] ), .B(n2100), .S0(n992), .Y(n1737) );
  CLKMX2X2 U1651 ( .A(\register[21][11] ), .B(n2105), .S0(n992), .Y(n1736) );
  CLKMX2X2 U1652 ( .A(\register[21][12] ), .B(n2110), .S0(n992), .Y(n1735) );
  CLKMX2X2 U1653 ( .A(\register[21][13] ), .B(n2115), .S0(n992), .Y(n1734) );
  CLKMX2X2 U1654 ( .A(\register[21][14] ), .B(n2120), .S0(n992), .Y(n1733) );
  CLKMX2X2 U1655 ( .A(\register[21][15] ), .B(n2125), .S0(n992), .Y(n1732) );
  CLKMX2X2 U1656 ( .A(\register[21][16] ), .B(n2130), .S0(n992), .Y(n1731) );
  CLKMX2X2 U1657 ( .A(\register[21][17] ), .B(n2135), .S0(n992), .Y(n1730) );
  CLKMX2X2 U1658 ( .A(\register[21][18] ), .B(n2140), .S0(n992), .Y(n1729) );
  CLKMX2X2 U1659 ( .A(\register[21][19] ), .B(n2145), .S0(n992), .Y(n1728) );
  CLKMX2X2 U1660 ( .A(\register[21][20] ), .B(n2150), .S0(n991), .Y(n1727) );
  CLKMX2X2 U1661 ( .A(\register[21][21] ), .B(n2155), .S0(n991), .Y(n1726) );
  CLKMX2X2 U1662 ( .A(\register[21][22] ), .B(n2160), .S0(n991), .Y(n1725) );
  CLKMX2X2 U1663 ( .A(\register[21][23] ), .B(n2165), .S0(n991), .Y(n1724) );
  CLKMX2X2 U1664 ( .A(\register[21][24] ), .B(n2170), .S0(n991), .Y(n1723) );
  CLKMX2X2 U1665 ( .A(\register[21][25] ), .B(n2175), .S0(n991), .Y(n1722) );
  CLKMX2X2 U1666 ( .A(\register[21][26] ), .B(n2180), .S0(n991), .Y(n1721) );
  CLKMX2X2 U1667 ( .A(\register[21][27] ), .B(n2185), .S0(n991), .Y(n1720) );
  CLKMX2X2 U1668 ( .A(\register[21][28] ), .B(n2190), .S0(n991), .Y(n1719) );
  CLKMX2X2 U1669 ( .A(\register[21][29] ), .B(n2195), .S0(n991), .Y(n1718) );
  CLKMX2X2 U1670 ( .A(\register[21][30] ), .B(n2200), .S0(n991), .Y(n1717) );
  CLKMX2X2 U1671 ( .A(\register[21][31] ), .B(n2205), .S0(n991), .Y(n1716) );
  CLKMX2X2 U1672 ( .A(\register[20][8] ), .B(n2090), .S0(n989), .Y(n1707) );
  CLKMX2X2 U1673 ( .A(\register[20][9] ), .B(n2095), .S0(n989), .Y(n1706) );
  CLKMX2X2 U1674 ( .A(\register[20][10] ), .B(n2100), .S0(n989), .Y(n1705) );
  CLKMX2X2 U1675 ( .A(\register[20][11] ), .B(n2105), .S0(n989), .Y(n1704) );
  CLKMX2X2 U1676 ( .A(\register[20][12] ), .B(n2110), .S0(n989), .Y(n1703) );
  CLKMX2X2 U1677 ( .A(\register[20][13] ), .B(n2115), .S0(n989), .Y(n1702) );
  CLKMX2X2 U1678 ( .A(\register[20][14] ), .B(n2120), .S0(n989), .Y(n1701) );
  CLKMX2X2 U1679 ( .A(\register[20][15] ), .B(n2125), .S0(n989), .Y(n1700) );
  CLKMX2X2 U1680 ( .A(\register[20][16] ), .B(n2130), .S0(n989), .Y(n1699) );
  CLKMX2X2 U1681 ( .A(\register[20][17] ), .B(n2135), .S0(n989), .Y(n1698) );
  CLKMX2X2 U1682 ( .A(\register[20][18] ), .B(n2140), .S0(n989), .Y(n1697) );
  CLKMX2X2 U1683 ( .A(\register[20][19] ), .B(n2145), .S0(n989), .Y(n1696) );
  CLKMX2X2 U1684 ( .A(\register[20][20] ), .B(n2150), .S0(n988), .Y(n1695) );
  CLKMX2X2 U1685 ( .A(\register[20][21] ), .B(n2155), .S0(n988), .Y(n1694) );
  CLKMX2X2 U1686 ( .A(\register[20][22] ), .B(n2160), .S0(n988), .Y(n1693) );
  CLKMX2X2 U1687 ( .A(\register[20][23] ), .B(n2165), .S0(n988), .Y(n1692) );
  CLKMX2X2 U1688 ( .A(\register[20][24] ), .B(n2170), .S0(n988), .Y(n1691) );
  CLKMX2X2 U1689 ( .A(\register[20][25] ), .B(n2175), .S0(n988), .Y(n1690) );
  CLKMX2X2 U1690 ( .A(\register[20][26] ), .B(n2180), .S0(n988), .Y(n1689) );
  CLKMX2X2 U1691 ( .A(\register[20][27] ), .B(n2185), .S0(n988), .Y(n1688) );
  CLKMX2X2 U1692 ( .A(\register[20][28] ), .B(n2190), .S0(n988), .Y(n1687) );
  CLKMX2X2 U1693 ( .A(\register[20][29] ), .B(n2195), .S0(n988), .Y(n1686) );
  CLKMX2X2 U1694 ( .A(\register[20][30] ), .B(n2200), .S0(n988), .Y(n1685) );
  CLKMX2X2 U1695 ( .A(\register[20][31] ), .B(n2205), .S0(n988), .Y(n1684) );
  CLKMX2X2 U1696 ( .A(\register[19][8] ), .B(n2091), .S0(n986), .Y(n1675) );
  CLKMX2X2 U1697 ( .A(\register[19][9] ), .B(n2096), .S0(n986), .Y(n1674) );
  CLKMX2X2 U1698 ( .A(\register[19][10] ), .B(n2101), .S0(n986), .Y(n1673) );
  CLKMX2X2 U1699 ( .A(\register[19][11] ), .B(n2106), .S0(n986), .Y(n1672) );
  CLKMX2X2 U1700 ( .A(\register[19][12] ), .B(n2111), .S0(n986), .Y(n1671) );
  CLKMX2X2 U1701 ( .A(\register[19][13] ), .B(n2116), .S0(n986), .Y(n1670) );
  CLKMX2X2 U1702 ( .A(\register[19][14] ), .B(n2121), .S0(n986), .Y(n1669) );
  CLKMX2X2 U1703 ( .A(\register[19][15] ), .B(n2126), .S0(n986), .Y(n1668) );
  CLKMX2X2 U1704 ( .A(\register[19][16] ), .B(n2131), .S0(n986), .Y(n1667) );
  CLKMX2X2 U1705 ( .A(\register[19][17] ), .B(n2136), .S0(n986), .Y(n1666) );
  CLKMX2X2 U1706 ( .A(\register[19][18] ), .B(n2141), .S0(n986), .Y(n1665) );
  CLKMX2X2 U1707 ( .A(\register[19][19] ), .B(n2146), .S0(n986), .Y(n1664) );
  CLKMX2X2 U1708 ( .A(\register[19][20] ), .B(n2151), .S0(n985), .Y(n1663) );
  CLKMX2X2 U1709 ( .A(\register[19][21] ), .B(n2156), .S0(n985), .Y(n1662) );
  CLKMX2X2 U1710 ( .A(\register[19][22] ), .B(n2161), .S0(n985), .Y(n1661) );
  CLKMX2X2 U1711 ( .A(\register[19][23] ), .B(n2166), .S0(n985), .Y(n1660) );
  CLKMX2X2 U1712 ( .A(\register[19][24] ), .B(n2171), .S0(n985), .Y(n1659) );
  CLKMX2X2 U1713 ( .A(\register[19][25] ), .B(n2176), .S0(n985), .Y(n1658) );
  CLKMX2X2 U1714 ( .A(\register[19][26] ), .B(n2181), .S0(n985), .Y(n1657) );
  CLKMX2X2 U1715 ( .A(\register[19][27] ), .B(n2186), .S0(n985), .Y(n1656) );
  CLKMX2X2 U1716 ( .A(\register[19][28] ), .B(n2191), .S0(n985), .Y(n1655) );
  CLKMX2X2 U1717 ( .A(\register[19][29] ), .B(n2196), .S0(n985), .Y(n1654) );
  CLKMX2X2 U1718 ( .A(\register[19][30] ), .B(n2201), .S0(n985), .Y(n1653) );
  CLKMX2X2 U1719 ( .A(\register[19][31] ), .B(n2205), .S0(n985), .Y(n1652) );
  CLKMX2X2 U1720 ( .A(\register[18][8] ), .B(n2091), .S0(n983), .Y(n1643) );
  CLKMX2X2 U1721 ( .A(\register[18][9] ), .B(n2096), .S0(n983), .Y(n1642) );
  CLKMX2X2 U1722 ( .A(\register[18][10] ), .B(n2101), .S0(n983), .Y(n1641) );
  CLKMX2X2 U1723 ( .A(\register[18][11] ), .B(n2106), .S0(n983), .Y(n1640) );
  CLKMX2X2 U1724 ( .A(\register[18][12] ), .B(n2111), .S0(n983), .Y(n1639) );
  CLKMX2X2 U1725 ( .A(\register[18][13] ), .B(n2116), .S0(n983), .Y(n1638) );
  CLKMX2X2 U1726 ( .A(\register[18][14] ), .B(n2121), .S0(n983), .Y(n1637) );
  CLKMX2X2 U1727 ( .A(\register[18][15] ), .B(n2126), .S0(n983), .Y(n1636) );
  CLKMX2X2 U1728 ( .A(\register[18][16] ), .B(n2131), .S0(n983), .Y(n1635) );
  CLKMX2X2 U1729 ( .A(\register[18][17] ), .B(n2136), .S0(n983), .Y(n1634) );
  CLKMX2X2 U1730 ( .A(\register[18][18] ), .B(n2141), .S0(n983), .Y(n1633) );
  CLKMX2X2 U1731 ( .A(\register[18][19] ), .B(n2146), .S0(n983), .Y(n1632) );
  CLKMX2X2 U1732 ( .A(\register[18][20] ), .B(n2151), .S0(n982), .Y(n1631) );
  CLKMX2X2 U1733 ( .A(\register[18][21] ), .B(n2156), .S0(n982), .Y(n1630) );
  CLKMX2X2 U1734 ( .A(\register[18][22] ), .B(n2161), .S0(n982), .Y(n1629) );
  CLKMX2X2 U1735 ( .A(\register[18][23] ), .B(n2166), .S0(n982), .Y(n1628) );
  CLKMX2X2 U1736 ( .A(\register[18][24] ), .B(n2171), .S0(n982), .Y(n1627) );
  CLKMX2X2 U1737 ( .A(\register[18][25] ), .B(n2176), .S0(n982), .Y(n1626) );
  CLKMX2X2 U1738 ( .A(\register[18][26] ), .B(n2181), .S0(n982), .Y(n1625) );
  CLKMX2X2 U1739 ( .A(\register[18][27] ), .B(n2186), .S0(n982), .Y(n1624) );
  CLKMX2X2 U1740 ( .A(\register[18][28] ), .B(n2191), .S0(n982), .Y(n1623) );
  CLKMX2X2 U1741 ( .A(\register[18][29] ), .B(n2196), .S0(n982), .Y(n1622) );
  CLKMX2X2 U1742 ( .A(\register[18][30] ), .B(n2201), .S0(n982), .Y(n1621) );
  CLKMX2X2 U1743 ( .A(\register[18][31] ), .B(n2205), .S0(n982), .Y(n1620) );
  CLKMX2X2 U1744 ( .A(\register[17][8] ), .B(n2091), .S0(n980), .Y(n1611) );
  CLKMX2X2 U1745 ( .A(\register[17][9] ), .B(n2096), .S0(n980), .Y(n1610) );
  CLKMX2X2 U1746 ( .A(\register[17][10] ), .B(n2101), .S0(n980), .Y(n1609) );
  CLKMX2X2 U1747 ( .A(\register[17][11] ), .B(n2106), .S0(n980), .Y(n1608) );
  CLKMX2X2 U1748 ( .A(\register[17][12] ), .B(n2111), .S0(n980), .Y(n1607) );
  CLKMX2X2 U1749 ( .A(\register[17][13] ), .B(n2116), .S0(n980), .Y(n1606) );
  CLKMX2X2 U1750 ( .A(\register[17][14] ), .B(n2121), .S0(n980), .Y(n1605) );
  CLKMX2X2 U1751 ( .A(\register[17][15] ), .B(n2126), .S0(n980), .Y(n1604) );
  CLKMX2X2 U1752 ( .A(\register[17][16] ), .B(n2131), .S0(n980), .Y(n1603) );
  CLKMX2X2 U1753 ( .A(\register[17][17] ), .B(n2136), .S0(n980), .Y(n1602) );
  CLKMX2X2 U1754 ( .A(\register[17][18] ), .B(n2141), .S0(n980), .Y(n1601) );
  CLKMX2X2 U1755 ( .A(\register[17][19] ), .B(n2146), .S0(n980), .Y(n1600) );
  CLKMX2X2 U1756 ( .A(\register[17][20] ), .B(n2151), .S0(n979), .Y(n1599) );
  CLKMX2X2 U1757 ( .A(\register[17][21] ), .B(n2156), .S0(n979), .Y(n1598) );
  CLKMX2X2 U1758 ( .A(\register[17][22] ), .B(n2161), .S0(n979), .Y(n1597) );
  CLKMX2X2 U1759 ( .A(\register[17][23] ), .B(n2166), .S0(n979), .Y(n1596) );
  CLKMX2X2 U1760 ( .A(\register[17][24] ), .B(n2171), .S0(n979), .Y(n1595) );
  CLKMX2X2 U1761 ( .A(\register[17][25] ), .B(n2176), .S0(n979), .Y(n1594) );
  CLKMX2X2 U1762 ( .A(\register[17][26] ), .B(n2181), .S0(n979), .Y(n1593) );
  CLKMX2X2 U1763 ( .A(\register[17][27] ), .B(n2186), .S0(n979), .Y(n1592) );
  CLKMX2X2 U1764 ( .A(\register[17][28] ), .B(n2191), .S0(n979), .Y(n1591) );
  CLKMX2X2 U1765 ( .A(\register[17][29] ), .B(n2196), .S0(n979), .Y(n1590) );
  CLKMX2X2 U1766 ( .A(\register[17][30] ), .B(n2201), .S0(n979), .Y(n1589) );
  CLKMX2X2 U1767 ( .A(\register[17][31] ), .B(n2205), .S0(n979), .Y(n1588) );
  CLKMX2X2 U1768 ( .A(\register[16][8] ), .B(n2091), .S0(n977), .Y(n1579) );
  CLKMX2X2 U1769 ( .A(\register[16][9] ), .B(n2096), .S0(n977), .Y(n1578) );
  CLKMX2X2 U1770 ( .A(\register[16][10] ), .B(n2101), .S0(n977), .Y(n1577) );
  CLKMX2X2 U1771 ( .A(\register[16][11] ), .B(n2106), .S0(n977), .Y(n1576) );
  CLKMX2X2 U1772 ( .A(\register[16][12] ), .B(n2111), .S0(n977), .Y(n1575) );
  CLKMX2X2 U1773 ( .A(\register[16][13] ), .B(n2116), .S0(n977), .Y(n1574) );
  CLKMX2X2 U1774 ( .A(\register[16][14] ), .B(n2121), .S0(n977), .Y(n1573) );
  CLKMX2X2 U1775 ( .A(\register[16][15] ), .B(n2126), .S0(n977), .Y(n1572) );
  CLKMX2X2 U1776 ( .A(\register[16][16] ), .B(n2131), .S0(n977), .Y(n1571) );
  CLKMX2X2 U1777 ( .A(\register[16][17] ), .B(n2136), .S0(n977), .Y(n1570) );
  CLKMX2X2 U1778 ( .A(\register[16][18] ), .B(n2141), .S0(n977), .Y(n1569) );
  CLKMX2X2 U1779 ( .A(\register[16][19] ), .B(n2146), .S0(n977), .Y(n1568) );
  CLKMX2X2 U1780 ( .A(\register[16][20] ), .B(n2151), .S0(n976), .Y(n1567) );
  CLKMX2X2 U1781 ( .A(\register[16][21] ), .B(n2156), .S0(n976), .Y(n1566) );
  CLKMX2X2 U1782 ( .A(\register[16][22] ), .B(n2161), .S0(n976), .Y(n1565) );
  CLKMX2X2 U1783 ( .A(\register[16][23] ), .B(n2166), .S0(n976), .Y(n1564) );
  CLKMX2X2 U1784 ( .A(\register[16][24] ), .B(n2171), .S0(n976), .Y(n1563) );
  CLKMX2X2 U1785 ( .A(\register[16][25] ), .B(n2176), .S0(n976), .Y(n1562) );
  CLKMX2X2 U1786 ( .A(\register[16][26] ), .B(n2181), .S0(n976), .Y(n1561) );
  CLKMX2X2 U1787 ( .A(\register[16][27] ), .B(n2186), .S0(n976), .Y(n1560) );
  CLKMX2X2 U1788 ( .A(\register[16][28] ), .B(n2191), .S0(n976), .Y(n1559) );
  CLKMX2X2 U1789 ( .A(\register[16][29] ), .B(n2196), .S0(n976), .Y(n1558) );
  CLKMX2X2 U1790 ( .A(\register[16][30] ), .B(n2201), .S0(n976), .Y(n1557) );
  CLKMX2X2 U1791 ( .A(\register[16][31] ), .B(n2205), .S0(n976), .Y(n1556) );
  CLKMX2X2 U1792 ( .A(\register[15][8] ), .B(n2091), .S0(n973), .Y(n1547) );
  CLKMX2X2 U1793 ( .A(\register[15][9] ), .B(n2096), .S0(n973), .Y(n1546) );
  CLKMX2X2 U1794 ( .A(\register[15][10] ), .B(n2101), .S0(n973), .Y(n1545) );
  CLKMX2X2 U1795 ( .A(\register[15][11] ), .B(n2106), .S0(n973), .Y(n1544) );
  CLKMX2X2 U1796 ( .A(\register[15][12] ), .B(n2111), .S0(n973), .Y(n1543) );
  CLKMX2X2 U1797 ( .A(\register[15][13] ), .B(n2116), .S0(n973), .Y(n1542) );
  CLKMX2X2 U1798 ( .A(\register[15][14] ), .B(n2121), .S0(n973), .Y(n1541) );
  CLKMX2X2 U1799 ( .A(\register[15][15] ), .B(n2126), .S0(n973), .Y(n1540) );
  CLKMX2X2 U1800 ( .A(\register[15][16] ), .B(n2131), .S0(n973), .Y(n1539) );
  CLKMX2X2 U1801 ( .A(\register[15][17] ), .B(n2136), .S0(n973), .Y(n1538) );
  CLKMX2X2 U1802 ( .A(\register[15][18] ), .B(n2141), .S0(n973), .Y(n1537) );
  CLKMX2X2 U1803 ( .A(\register[15][19] ), .B(n2146), .S0(n973), .Y(n1536) );
  CLKMX2X2 U1804 ( .A(\register[15][20] ), .B(n2151), .S0(n972), .Y(n1535) );
  CLKMX2X2 U1805 ( .A(\register[15][21] ), .B(n2156), .S0(n972), .Y(n1534) );
  CLKMX2X2 U1806 ( .A(\register[15][22] ), .B(n2161), .S0(n972), .Y(n1533) );
  CLKMX2X2 U1807 ( .A(\register[15][23] ), .B(n2166), .S0(n972), .Y(n1532) );
  CLKMX2X2 U1808 ( .A(\register[15][24] ), .B(n2171), .S0(n972), .Y(n1531) );
  CLKMX2X2 U1809 ( .A(\register[15][25] ), .B(n2176), .S0(n972), .Y(n1530) );
  CLKMX2X2 U1810 ( .A(\register[15][26] ), .B(n2181), .S0(n972), .Y(n1529) );
  CLKMX2X2 U1811 ( .A(\register[15][27] ), .B(n2186), .S0(n972), .Y(n1528) );
  CLKMX2X2 U1812 ( .A(\register[15][28] ), .B(n2191), .S0(n972), .Y(n1527) );
  CLKMX2X2 U1813 ( .A(\register[15][29] ), .B(n2196), .S0(n972), .Y(n1526) );
  CLKMX2X2 U1814 ( .A(\register[15][30] ), .B(n2201), .S0(n972), .Y(n1525) );
  CLKMX2X2 U1815 ( .A(\register[15][31] ), .B(n2205), .S0(n972), .Y(n1524) );
  CLKMX2X2 U1816 ( .A(\register[14][8] ), .B(n2091), .S0(n970), .Y(n1515) );
  CLKMX2X2 U1817 ( .A(\register[14][9] ), .B(n2096), .S0(n970), .Y(n1514) );
  CLKMX2X2 U1818 ( .A(\register[14][10] ), .B(n2101), .S0(n970), .Y(n1513) );
  CLKMX2X2 U1819 ( .A(\register[14][11] ), .B(n2106), .S0(n970), .Y(n1512) );
  CLKMX2X2 U1820 ( .A(\register[14][12] ), .B(n2111), .S0(n970), .Y(n1511) );
  CLKMX2X2 U1821 ( .A(\register[14][13] ), .B(n2116), .S0(n970), .Y(n1510) );
  CLKMX2X2 U1822 ( .A(\register[14][14] ), .B(n2121), .S0(n970), .Y(n1509) );
  CLKMX2X2 U1823 ( .A(\register[14][15] ), .B(n2126), .S0(n970), .Y(n1508) );
  CLKMX2X2 U1824 ( .A(\register[14][16] ), .B(n2131), .S0(n970), .Y(n1507) );
  CLKMX2X2 U1825 ( .A(\register[14][17] ), .B(n2136), .S0(n970), .Y(n1506) );
  CLKMX2X2 U1826 ( .A(\register[14][18] ), .B(n2141), .S0(n970), .Y(n1505) );
  CLKMX2X2 U1827 ( .A(\register[14][19] ), .B(n2146), .S0(n970), .Y(n1504) );
  CLKMX2X2 U1828 ( .A(\register[14][20] ), .B(n2151), .S0(n969), .Y(n1503) );
  CLKMX2X2 U1829 ( .A(\register[14][21] ), .B(n2156), .S0(n969), .Y(n1502) );
  CLKMX2X2 U1830 ( .A(\register[14][22] ), .B(n2161), .S0(n969), .Y(n1501) );
  CLKMX2X2 U1831 ( .A(\register[14][23] ), .B(n2166), .S0(n969), .Y(n1500) );
  CLKMX2X2 U1832 ( .A(\register[14][24] ), .B(n2171), .S0(n969), .Y(n1499) );
  CLKMX2X2 U1833 ( .A(\register[14][25] ), .B(n2176), .S0(n969), .Y(n1498) );
  CLKMX2X2 U1834 ( .A(\register[14][26] ), .B(n2181), .S0(n969), .Y(n1497) );
  CLKMX2X2 U1835 ( .A(\register[14][27] ), .B(n2186), .S0(n969), .Y(n1496) );
  CLKMX2X2 U1836 ( .A(\register[14][28] ), .B(n2191), .S0(n969), .Y(n1495) );
  CLKMX2X2 U1837 ( .A(\register[14][29] ), .B(n2196), .S0(n969), .Y(n1494) );
  CLKMX2X2 U1838 ( .A(\register[14][30] ), .B(n2201), .S0(n969), .Y(n1493) );
  CLKMX2X2 U1839 ( .A(\register[14][31] ), .B(n2205), .S0(n969), .Y(n1492) );
  CLKMX2X2 U1840 ( .A(\register[13][8] ), .B(n2091), .S0(n967), .Y(n1483) );
  CLKMX2X2 U1841 ( .A(\register[13][9] ), .B(n2096), .S0(n967), .Y(n1482) );
  CLKMX2X2 U1842 ( .A(\register[13][10] ), .B(n2101), .S0(n967), .Y(n1481) );
  CLKMX2X2 U1843 ( .A(\register[13][11] ), .B(n2106), .S0(n967), .Y(n1480) );
  CLKMX2X2 U1844 ( .A(\register[13][12] ), .B(n2111), .S0(n967), .Y(n1479) );
  CLKMX2X2 U1845 ( .A(\register[13][13] ), .B(n2116), .S0(n967), .Y(n1478) );
  CLKMX2X2 U1846 ( .A(\register[13][14] ), .B(n2121), .S0(n967), .Y(n1477) );
  CLKMX2X2 U1847 ( .A(\register[13][15] ), .B(n2126), .S0(n967), .Y(n1476) );
  CLKMX2X2 U1848 ( .A(\register[13][16] ), .B(n2131), .S0(n967), .Y(n1475) );
  CLKMX2X2 U1849 ( .A(\register[13][17] ), .B(n2136), .S0(n967), .Y(n1474) );
  CLKMX2X2 U1850 ( .A(\register[13][18] ), .B(n2141), .S0(n967), .Y(n1473) );
  CLKMX2X2 U1851 ( .A(\register[13][19] ), .B(n2146), .S0(n967), .Y(n1472) );
  CLKMX2X2 U1852 ( .A(\register[13][20] ), .B(n2151), .S0(n966), .Y(n1471) );
  CLKMX2X2 U1853 ( .A(\register[13][21] ), .B(n2156), .S0(n966), .Y(n1470) );
  CLKMX2X2 U1854 ( .A(\register[13][22] ), .B(n2161), .S0(n966), .Y(n1469) );
  CLKMX2X2 U1855 ( .A(\register[13][23] ), .B(n2166), .S0(n966), .Y(n1468) );
  CLKMX2X2 U1856 ( .A(\register[13][24] ), .B(n2171), .S0(n966), .Y(n1467) );
  CLKMX2X2 U1857 ( .A(\register[13][25] ), .B(n2176), .S0(n966), .Y(n1466) );
  CLKMX2X2 U1858 ( .A(\register[13][26] ), .B(n2181), .S0(n966), .Y(n1465) );
  CLKMX2X2 U1859 ( .A(\register[13][27] ), .B(n2186), .S0(n966), .Y(n1464) );
  CLKMX2X2 U1860 ( .A(\register[13][28] ), .B(n2191), .S0(n966), .Y(n1463) );
  CLKMX2X2 U1861 ( .A(\register[13][29] ), .B(n2196), .S0(n966), .Y(n1462) );
  CLKMX2X2 U1862 ( .A(\register[13][30] ), .B(n2201), .S0(n966), .Y(n1461) );
  CLKMX2X2 U1863 ( .A(\register[13][31] ), .B(n2205), .S0(n966), .Y(n1460) );
  CLKMX2X2 U1864 ( .A(\register[12][8] ), .B(n2091), .S0(n964), .Y(n1451) );
  CLKMX2X2 U1865 ( .A(\register[12][9] ), .B(n2096), .S0(n964), .Y(n1450) );
  CLKMX2X2 U1866 ( .A(\register[12][10] ), .B(n2101), .S0(n964), .Y(n1449) );
  CLKMX2X2 U1867 ( .A(\register[12][11] ), .B(n2106), .S0(n964), .Y(n1448) );
  CLKMX2X2 U1868 ( .A(\register[12][12] ), .B(n2111), .S0(n964), .Y(n1447) );
  CLKMX2X2 U1869 ( .A(\register[12][13] ), .B(n2116), .S0(n964), .Y(n1446) );
  CLKMX2X2 U1870 ( .A(\register[12][14] ), .B(n2121), .S0(n964), .Y(n1445) );
  CLKMX2X2 U1871 ( .A(\register[12][15] ), .B(n2126), .S0(n964), .Y(n1444) );
  CLKMX2X2 U1872 ( .A(\register[12][16] ), .B(n2131), .S0(n964), .Y(n1443) );
  CLKMX2X2 U1873 ( .A(\register[12][17] ), .B(n2136), .S0(n964), .Y(n1442) );
  CLKMX2X2 U1874 ( .A(\register[12][18] ), .B(n2141), .S0(n964), .Y(n1441) );
  CLKMX2X2 U1875 ( .A(\register[12][19] ), .B(n2146), .S0(n964), .Y(n1440) );
  CLKMX2X2 U1876 ( .A(\register[12][20] ), .B(n2151), .S0(n963), .Y(n1439) );
  CLKMX2X2 U1877 ( .A(\register[12][21] ), .B(n2156), .S0(n963), .Y(n1438) );
  CLKMX2X2 U1878 ( .A(\register[12][22] ), .B(n2161), .S0(n963), .Y(n1437) );
  CLKMX2X2 U1879 ( .A(\register[12][23] ), .B(n2166), .S0(n963), .Y(n1436) );
  CLKMX2X2 U1880 ( .A(\register[12][24] ), .B(n2171), .S0(n963), .Y(n1435) );
  CLKMX2X2 U1881 ( .A(\register[12][25] ), .B(n2176), .S0(n963), .Y(n1434) );
  CLKMX2X2 U1882 ( .A(\register[12][26] ), .B(n2181), .S0(n963), .Y(n1433) );
  CLKMX2X2 U1883 ( .A(\register[12][27] ), .B(n2186), .S0(n963), .Y(n1432) );
  CLKMX2X2 U1884 ( .A(\register[12][28] ), .B(n2191), .S0(n963), .Y(n1431) );
  CLKMX2X2 U1885 ( .A(\register[12][29] ), .B(n2196), .S0(n963), .Y(n1430) );
  CLKMX2X2 U1886 ( .A(\register[12][30] ), .B(n2201), .S0(n963), .Y(n1429) );
  CLKMX2X2 U1887 ( .A(\register[12][31] ), .B(n2205), .S0(n963), .Y(n1428) );
  CLKMX2X2 U1888 ( .A(\register[11][8] ), .B(n2091), .S0(n961), .Y(n1419) );
  CLKMX2X2 U1889 ( .A(\register[11][9] ), .B(n2096), .S0(n961), .Y(n1418) );
  CLKMX2X2 U1890 ( .A(\register[11][10] ), .B(n2101), .S0(n961), .Y(n1417) );
  CLKMX2X2 U1891 ( .A(\register[11][11] ), .B(n2106), .S0(n961), .Y(n1416) );
  CLKMX2X2 U1892 ( .A(\register[11][12] ), .B(n2111), .S0(n961), .Y(n1415) );
  CLKMX2X2 U1893 ( .A(\register[11][13] ), .B(n2116), .S0(n961), .Y(n1414) );
  CLKMX2X2 U1894 ( .A(\register[11][14] ), .B(n2121), .S0(n961), .Y(n1413) );
  CLKMX2X2 U1895 ( .A(\register[11][15] ), .B(n2126), .S0(n961), .Y(n1412) );
  CLKMX2X2 U1896 ( .A(\register[11][16] ), .B(n2131), .S0(n961), .Y(n1411) );
  CLKMX2X2 U1897 ( .A(\register[11][17] ), .B(n2136), .S0(n961), .Y(n1410) );
  CLKMX2X2 U1898 ( .A(\register[11][18] ), .B(n2141), .S0(n961), .Y(n1409) );
  CLKMX2X2 U1899 ( .A(\register[11][19] ), .B(n2146), .S0(n961), .Y(n1408) );
  CLKMX2X2 U1900 ( .A(\register[11][20] ), .B(n2151), .S0(n960), .Y(n1407) );
  CLKMX2X2 U1901 ( .A(\register[11][21] ), .B(n2156), .S0(n960), .Y(n1406) );
  CLKMX2X2 U1902 ( .A(\register[11][22] ), .B(n2161), .S0(n960), .Y(n1405) );
  CLKMX2X2 U1903 ( .A(\register[11][23] ), .B(n2166), .S0(n960), .Y(n1404) );
  CLKMX2X2 U1904 ( .A(\register[11][24] ), .B(n2171), .S0(n960), .Y(n1403) );
  CLKMX2X2 U1905 ( .A(\register[11][25] ), .B(n2176), .S0(n960), .Y(n1402) );
  CLKMX2X2 U1906 ( .A(\register[11][26] ), .B(n2181), .S0(n960), .Y(n1401) );
  CLKMX2X2 U1907 ( .A(\register[11][27] ), .B(n2186), .S0(n960), .Y(n1400) );
  CLKMX2X2 U1908 ( .A(\register[11][28] ), .B(n2191), .S0(n960), .Y(n1399) );
  CLKMX2X2 U1909 ( .A(\register[11][29] ), .B(n2196), .S0(n960), .Y(n1398) );
  CLKMX2X2 U1910 ( .A(\register[11][30] ), .B(n2201), .S0(n960), .Y(n1397) );
  CLKMX2X2 U1911 ( .A(\register[11][31] ), .B(n2205), .S0(n960), .Y(n1396) );
  CLKMX2X2 U1912 ( .A(\register[10][8] ), .B(n2091), .S0(n958), .Y(n1387) );
  CLKMX2X2 U1913 ( .A(\register[10][9] ), .B(n2096), .S0(n958), .Y(n1386) );
  CLKMX2X2 U1914 ( .A(\register[10][10] ), .B(n2101), .S0(n958), .Y(n1385) );
  CLKMX2X2 U1915 ( .A(\register[10][11] ), .B(n2106), .S0(n958), .Y(n1384) );
  CLKMX2X2 U1916 ( .A(\register[10][12] ), .B(n2111), .S0(n958), .Y(n1383) );
  CLKMX2X2 U1917 ( .A(\register[10][13] ), .B(n2116), .S0(n958), .Y(n1382) );
  CLKMX2X2 U1918 ( .A(\register[10][14] ), .B(n2121), .S0(n958), .Y(n1381) );
  CLKMX2X2 U1919 ( .A(\register[10][15] ), .B(n2126), .S0(n958), .Y(n1380) );
  CLKMX2X2 U1920 ( .A(\register[10][16] ), .B(n2131), .S0(n958), .Y(n1379) );
  CLKMX2X2 U1921 ( .A(\register[10][17] ), .B(n2136), .S0(n958), .Y(n1378) );
  CLKMX2X2 U1922 ( .A(\register[10][18] ), .B(n2141), .S0(n958), .Y(n1377) );
  CLKMX2X2 U1923 ( .A(\register[10][19] ), .B(n2146), .S0(n958), .Y(n1376) );
  CLKMX2X2 U1924 ( .A(\register[10][20] ), .B(n2151), .S0(n957), .Y(n1375) );
  CLKMX2X2 U1925 ( .A(\register[10][21] ), .B(n2156), .S0(n957), .Y(n1374) );
  CLKMX2X2 U1926 ( .A(\register[10][22] ), .B(n2161), .S0(n957), .Y(n1373) );
  CLKMX2X2 U1927 ( .A(\register[10][23] ), .B(n2166), .S0(n957), .Y(n1372) );
  CLKMX2X2 U1928 ( .A(\register[10][24] ), .B(n2171), .S0(n957), .Y(n1371) );
  CLKMX2X2 U1929 ( .A(\register[10][25] ), .B(n2176), .S0(n957), .Y(n1370) );
  CLKMX2X2 U1930 ( .A(\register[10][26] ), .B(n2181), .S0(n957), .Y(n1369) );
  CLKMX2X2 U1931 ( .A(\register[10][27] ), .B(n2186), .S0(n957), .Y(n1368) );
  CLKMX2X2 U1932 ( .A(\register[10][28] ), .B(n2191), .S0(n957), .Y(n1367) );
  CLKMX2X2 U1933 ( .A(\register[10][29] ), .B(n2196), .S0(n957), .Y(n1366) );
  CLKMX2X2 U1934 ( .A(\register[10][30] ), .B(n2201), .S0(n957), .Y(n1365) );
  CLKMX2X2 U1935 ( .A(\register[10][31] ), .B(n2205), .S0(n957), .Y(n1364) );
  CLKMX2X2 U1936 ( .A(\register[9][8] ), .B(n2091), .S0(n955), .Y(n1355) );
  CLKMX2X2 U1937 ( .A(\register[9][9] ), .B(n2096), .S0(n955), .Y(n1354) );
  CLKMX2X2 U1938 ( .A(\register[9][10] ), .B(n2101), .S0(n955), .Y(n1353) );
  CLKMX2X2 U1939 ( .A(\register[9][11] ), .B(n2106), .S0(n955), .Y(n1352) );
  CLKMX2X2 U1940 ( .A(\register[9][12] ), .B(n2111), .S0(n955), .Y(n1351) );
  CLKMX2X2 U1941 ( .A(\register[9][13] ), .B(n2116), .S0(n955), .Y(n1350) );
  CLKMX2X2 U1942 ( .A(\register[9][14] ), .B(n2121), .S0(n955), .Y(n1349) );
  CLKMX2X2 U1943 ( .A(\register[9][15] ), .B(n2126), .S0(n955), .Y(n1348) );
  CLKMX2X2 U1944 ( .A(\register[9][16] ), .B(n2131), .S0(n955), .Y(n1347) );
  CLKMX2X2 U1945 ( .A(\register[9][17] ), .B(n2136), .S0(n955), .Y(n1346) );
  CLKMX2X2 U1946 ( .A(\register[9][18] ), .B(n2141), .S0(n955), .Y(n1345) );
  CLKMX2X2 U1947 ( .A(\register[9][19] ), .B(n2146), .S0(n955), .Y(n1344) );
  CLKMX2X2 U1948 ( .A(\register[9][20] ), .B(n2151), .S0(n954), .Y(n1343) );
  CLKMX2X2 U1949 ( .A(\register[9][21] ), .B(n2156), .S0(n954), .Y(n1342) );
  CLKMX2X2 U1950 ( .A(\register[9][22] ), .B(n2161), .S0(n954), .Y(n1341) );
  CLKMX2X2 U1951 ( .A(\register[9][23] ), .B(n2166), .S0(n954), .Y(n1340) );
  CLKMX2X2 U1952 ( .A(\register[9][24] ), .B(n2171), .S0(n954), .Y(n1339) );
  CLKMX2X2 U1953 ( .A(\register[9][25] ), .B(n2176), .S0(n954), .Y(n1338) );
  CLKMX2X2 U1954 ( .A(\register[9][26] ), .B(n2181), .S0(n954), .Y(n1337) );
  CLKMX2X2 U1955 ( .A(\register[9][27] ), .B(n2186), .S0(n954), .Y(n1336) );
  CLKMX2X2 U1956 ( .A(\register[9][28] ), .B(n2191), .S0(n954), .Y(n1335) );
  CLKMX2X2 U1957 ( .A(\register[9][29] ), .B(n2196), .S0(n954), .Y(n1334) );
  CLKMX2X2 U1958 ( .A(\register[9][30] ), .B(n2201), .S0(n954), .Y(n1333) );
  CLKMX2X2 U1959 ( .A(\register[9][31] ), .B(n2205), .S0(n954), .Y(n1332) );
  CLKMX2X2 U1960 ( .A(\register[8][8] ), .B(n2091), .S0(n952), .Y(n1323) );
  CLKMX2X2 U1961 ( .A(\register[8][9] ), .B(n2096), .S0(n952), .Y(n1322) );
  CLKMX2X2 U1962 ( .A(\register[8][10] ), .B(n2101), .S0(n952), .Y(n1321) );
  CLKMX2X2 U1963 ( .A(\register[8][11] ), .B(n2106), .S0(n952), .Y(n1320) );
  CLKMX2X2 U1964 ( .A(\register[8][12] ), .B(n2111), .S0(n952), .Y(n1319) );
  CLKMX2X2 U1965 ( .A(\register[8][13] ), .B(n2116), .S0(n952), .Y(n1318) );
  CLKMX2X2 U1966 ( .A(\register[8][14] ), .B(n2121), .S0(n952), .Y(n1317) );
  CLKMX2X2 U1967 ( .A(\register[8][15] ), .B(n2126), .S0(n952), .Y(n1316) );
  CLKMX2X2 U1968 ( .A(\register[8][16] ), .B(n2131), .S0(n952), .Y(n1315) );
  CLKMX2X2 U1969 ( .A(\register[8][17] ), .B(n2136), .S0(n952), .Y(n1314) );
  CLKMX2X2 U1970 ( .A(\register[8][18] ), .B(n2141), .S0(n952), .Y(n1313) );
  CLKMX2X2 U1971 ( .A(\register[8][19] ), .B(n2146), .S0(n952), .Y(n1312) );
  CLKMX2X2 U1972 ( .A(\register[8][20] ), .B(n2151), .S0(n951), .Y(n1311) );
  CLKMX2X2 U1973 ( .A(\register[8][21] ), .B(n2156), .S0(n951), .Y(n1310) );
  CLKMX2X2 U1974 ( .A(\register[8][22] ), .B(n2161), .S0(n951), .Y(n1309) );
  CLKMX2X2 U1975 ( .A(\register[8][23] ), .B(n2166), .S0(n951), .Y(n1308) );
  CLKMX2X2 U1976 ( .A(\register[8][24] ), .B(n2171), .S0(n951), .Y(n1307) );
  CLKMX2X2 U1977 ( .A(\register[8][25] ), .B(n2176), .S0(n951), .Y(n1306) );
  CLKMX2X2 U1978 ( .A(\register[8][26] ), .B(n2181), .S0(n951), .Y(n1305) );
  CLKMX2X2 U1979 ( .A(\register[8][27] ), .B(n2186), .S0(n951), .Y(n1304) );
  CLKMX2X2 U1980 ( .A(\register[8][28] ), .B(n2191), .S0(n951), .Y(n1303) );
  CLKMX2X2 U1981 ( .A(\register[8][29] ), .B(n2196), .S0(n951), .Y(n1302) );
  CLKMX2X2 U1982 ( .A(\register[8][30] ), .B(n2201), .S0(n951), .Y(n1301) );
  CLKMX2X2 U1983 ( .A(\register[8][31] ), .B(n2205), .S0(n951), .Y(n1300) );
  CLKMX2X2 U1984 ( .A(\register[7][8] ), .B(n2092), .S0(n949), .Y(n1291) );
  CLKMX2X2 U1985 ( .A(\register[7][9] ), .B(n2097), .S0(n949), .Y(n1290) );
  CLKMX2X2 U1986 ( .A(\register[7][10] ), .B(n2102), .S0(n949), .Y(n1289) );
  CLKMX2X2 U1987 ( .A(\register[7][11] ), .B(n2107), .S0(n949), .Y(n1288) );
  CLKMX2X2 U1988 ( .A(\register[7][12] ), .B(n2112), .S0(n949), .Y(n1287) );
  CLKMX2X2 U1989 ( .A(\register[7][13] ), .B(n2117), .S0(n949), .Y(n1286) );
  CLKMX2X2 U1990 ( .A(\register[7][14] ), .B(n2122), .S0(n949), .Y(n1285) );
  CLKMX2X2 U1991 ( .A(\register[7][15] ), .B(n2127), .S0(n949), .Y(n1284) );
  CLKMX2X2 U1992 ( .A(\register[7][16] ), .B(n2132), .S0(n949), .Y(n1283) );
  CLKMX2X2 U1993 ( .A(\register[7][17] ), .B(n2137), .S0(n949), .Y(n1282) );
  CLKMX2X2 U1994 ( .A(\register[7][18] ), .B(n2142), .S0(n949), .Y(n1281) );
  CLKMX2X2 U1995 ( .A(\register[7][19] ), .B(n2147), .S0(n949), .Y(n1280) );
  CLKMX2X2 U1996 ( .A(\register[7][20] ), .B(n2152), .S0(n948), .Y(n1279) );
  CLKMX2X2 U1997 ( .A(\register[7][21] ), .B(n2157), .S0(n948), .Y(n1278) );
  CLKMX2X2 U1998 ( .A(\register[7][22] ), .B(n2162), .S0(n948), .Y(n1277) );
  CLKMX2X2 U1999 ( .A(\register[7][23] ), .B(n2167), .S0(n948), .Y(n1276) );
  CLKMX2X2 U2000 ( .A(\register[7][24] ), .B(n2172), .S0(n948), .Y(n1275) );
  CLKMX2X2 U2001 ( .A(\register[7][25] ), .B(n2177), .S0(n948), .Y(n1274) );
  CLKMX2X2 U2002 ( .A(\register[7][26] ), .B(n2182), .S0(n948), .Y(n1273) );
  CLKMX2X2 U2003 ( .A(\register[7][27] ), .B(n2187), .S0(n948), .Y(n1272) );
  CLKMX2X2 U2004 ( .A(\register[7][28] ), .B(n2192), .S0(n948), .Y(n1271) );
  CLKMX2X2 U2005 ( .A(\register[7][29] ), .B(n2197), .S0(n948), .Y(n1270) );
  CLKMX2X2 U2006 ( .A(\register[7][30] ), .B(n2202), .S0(n948), .Y(n1269) );
  CLKMX2X2 U2007 ( .A(\register[7][31] ), .B(n2205), .S0(n948), .Y(n1268) );
  CLKMX2X2 U2008 ( .A(\register[6][8] ), .B(n2092), .S0(n946), .Y(n1259) );
  CLKMX2X2 U2009 ( .A(\register[6][9] ), .B(n2097), .S0(n946), .Y(n1258) );
  CLKMX2X2 U2010 ( .A(\register[6][10] ), .B(n2102), .S0(n946), .Y(n1257) );
  CLKMX2X2 U2011 ( .A(\register[6][11] ), .B(n2107), .S0(n946), .Y(n1256) );
  CLKMX2X2 U2012 ( .A(\register[6][12] ), .B(n2112), .S0(n946), .Y(n1255) );
  CLKMX2X2 U2013 ( .A(\register[6][13] ), .B(n2117), .S0(n946), .Y(n1254) );
  CLKMX2X2 U2014 ( .A(\register[6][14] ), .B(n2122), .S0(n946), .Y(n1253) );
  CLKMX2X2 U2015 ( .A(\register[6][15] ), .B(n2127), .S0(n946), .Y(n1252) );
  CLKMX2X2 U2016 ( .A(\register[6][16] ), .B(n2132), .S0(n946), .Y(n1251) );
  CLKMX2X2 U2017 ( .A(\register[6][17] ), .B(n2137), .S0(n946), .Y(n1250) );
  CLKMX2X2 U2018 ( .A(\register[6][18] ), .B(n2142), .S0(n946), .Y(n1249) );
  CLKMX2X2 U2019 ( .A(\register[6][19] ), .B(n2147), .S0(n946), .Y(n1248) );
  CLKMX2X2 U2020 ( .A(\register[6][20] ), .B(n2152), .S0(n945), .Y(n1247) );
  CLKMX2X2 U2021 ( .A(\register[6][21] ), .B(n2157), .S0(n945), .Y(n1246) );
  CLKMX2X2 U2022 ( .A(\register[6][22] ), .B(n2162), .S0(n945), .Y(n1245) );
  CLKMX2X2 U2023 ( .A(\register[6][23] ), .B(n2167), .S0(n945), .Y(n1244) );
  CLKMX2X2 U2024 ( .A(\register[6][24] ), .B(n2172), .S0(n945), .Y(n1243) );
  CLKMX2X2 U2025 ( .A(\register[6][25] ), .B(n2177), .S0(n945), .Y(n1242) );
  CLKMX2X2 U2026 ( .A(\register[6][26] ), .B(n2182), .S0(n945), .Y(n1241) );
  CLKMX2X2 U2027 ( .A(\register[6][27] ), .B(n2187), .S0(n945), .Y(n1240) );
  CLKMX2X2 U2028 ( .A(\register[6][28] ), .B(n2192), .S0(n945), .Y(n1239) );
  CLKMX2X2 U2029 ( .A(\register[6][29] ), .B(n2197), .S0(n945), .Y(n1238) );
  CLKMX2X2 U2030 ( .A(\register[6][30] ), .B(n2202), .S0(n945), .Y(n1237) );
  CLKMX2X2 U2031 ( .A(\register[6][31] ), .B(n2205), .S0(n945), .Y(n1236) );
  CLKMX2X2 U2032 ( .A(\register[5][8] ), .B(n2092), .S0(n943), .Y(n1227) );
  CLKMX2X2 U2033 ( .A(\register[5][9] ), .B(n2097), .S0(n943), .Y(n1226) );
  CLKMX2X2 U2034 ( .A(\register[5][10] ), .B(n2102), .S0(n943), .Y(n1225) );
  CLKMX2X2 U2035 ( .A(\register[5][11] ), .B(n2107), .S0(n943), .Y(n1224) );
  CLKMX2X2 U2036 ( .A(\register[5][12] ), .B(n2112), .S0(n943), .Y(n1223) );
  CLKMX2X2 U2037 ( .A(\register[5][13] ), .B(n2117), .S0(n943), .Y(n1222) );
  CLKMX2X2 U2038 ( .A(\register[5][14] ), .B(n2122), .S0(n943), .Y(n1221) );
  CLKMX2X2 U2039 ( .A(\register[5][15] ), .B(n2127), .S0(n943), .Y(n1220) );
  CLKMX2X2 U2040 ( .A(\register[5][16] ), .B(n2132), .S0(n943), .Y(n1219) );
  CLKMX2X2 U2041 ( .A(\register[5][17] ), .B(n2137), .S0(n943), .Y(n1218) );
  CLKMX2X2 U2042 ( .A(\register[5][18] ), .B(n2142), .S0(n943), .Y(n1217) );
  CLKMX2X2 U2043 ( .A(\register[5][19] ), .B(n2147), .S0(n943), .Y(n1216) );
  CLKMX2X2 U2044 ( .A(\register[5][20] ), .B(n2152), .S0(n942), .Y(n1215) );
  CLKMX2X2 U2045 ( .A(\register[5][21] ), .B(n2157), .S0(n942), .Y(n1214) );
  CLKMX2X2 U2046 ( .A(\register[5][22] ), .B(n2162), .S0(n942), .Y(n1213) );
  CLKMX2X2 U2047 ( .A(\register[5][23] ), .B(n2167), .S0(n942), .Y(n1212) );
  CLKMX2X2 U2048 ( .A(\register[5][24] ), .B(n2172), .S0(n942), .Y(n1211) );
  CLKMX2X2 U2049 ( .A(\register[5][25] ), .B(n2177), .S0(n942), .Y(n1210) );
  CLKMX2X2 U2050 ( .A(\register[5][26] ), .B(n2182), .S0(n942), .Y(n1209) );
  CLKMX2X2 U2051 ( .A(\register[5][27] ), .B(n2187), .S0(n942), .Y(n1208) );
  CLKMX2X2 U2052 ( .A(\register[5][28] ), .B(n2192), .S0(n942), .Y(n1207) );
  CLKMX2X2 U2053 ( .A(\register[5][29] ), .B(n2197), .S0(n942), .Y(n1206) );
  CLKMX2X2 U2054 ( .A(\register[5][30] ), .B(n2202), .S0(n942), .Y(n1205) );
  CLKMX2X2 U2055 ( .A(\register[5][31] ), .B(n2205), .S0(n942), .Y(n1204) );
  CLKMX2X2 U2056 ( .A(\register[4][8] ), .B(n2092), .S0(n939), .Y(n1195) );
  CLKMX2X2 U2057 ( .A(\register[4][9] ), .B(n2097), .S0(n939), .Y(n1194) );
  CLKMX2X2 U2058 ( .A(\register[4][10] ), .B(n2102), .S0(n939), .Y(n1193) );
  CLKMX2X2 U2059 ( .A(\register[4][11] ), .B(n2107), .S0(n939), .Y(n1192) );
  CLKMX2X2 U2060 ( .A(\register[4][12] ), .B(n2112), .S0(n939), .Y(n1191) );
  CLKMX2X2 U2061 ( .A(\register[4][13] ), .B(n2117), .S0(n939), .Y(n1190) );
  CLKMX2X2 U2062 ( .A(\register[4][14] ), .B(n2122), .S0(n939), .Y(n1189) );
  CLKMX2X2 U2063 ( .A(\register[4][15] ), .B(n2127), .S0(n939), .Y(n1188) );
  CLKMX2X2 U2064 ( .A(\register[4][16] ), .B(n2132), .S0(n939), .Y(n1187) );
  CLKMX2X2 U2065 ( .A(\register[4][17] ), .B(n2137), .S0(n939), .Y(n1186) );
  CLKMX2X2 U2066 ( .A(\register[4][18] ), .B(n2142), .S0(n939), .Y(n1185) );
  CLKMX2X2 U2067 ( .A(\register[4][19] ), .B(n2147), .S0(n939), .Y(n1184) );
  CLKMX2X2 U2068 ( .A(\register[4][20] ), .B(n2152), .S0(n938), .Y(n1183) );
  CLKMX2X2 U2069 ( .A(\register[4][21] ), .B(n2157), .S0(n938), .Y(n1182) );
  CLKMX2X2 U2070 ( .A(\register[4][22] ), .B(n2162), .S0(n938), .Y(n1181) );
  CLKMX2X2 U2071 ( .A(\register[4][23] ), .B(n2167), .S0(n938), .Y(n1180) );
  CLKMX2X2 U2072 ( .A(\register[4][24] ), .B(n2172), .S0(n938), .Y(n1179) );
  CLKMX2X2 U2073 ( .A(\register[4][25] ), .B(n2177), .S0(n938), .Y(n1178) );
  CLKMX2X2 U2074 ( .A(\register[4][26] ), .B(n2182), .S0(n938), .Y(n1177) );
  CLKMX2X2 U2075 ( .A(\register[4][27] ), .B(n2187), .S0(n938), .Y(n1176) );
  CLKMX2X2 U2076 ( .A(\register[4][28] ), .B(n2192), .S0(n938), .Y(n1175) );
  CLKMX2X2 U2077 ( .A(\register[4][29] ), .B(n2197), .S0(n938), .Y(n1174) );
  CLKMX2X2 U2078 ( .A(\register[4][30] ), .B(n2202), .S0(n938), .Y(n1173) );
  CLKMX2X2 U2079 ( .A(\register[4][31] ), .B(n2205), .S0(n938), .Y(n1172) );
  CLKMX2X2 U2080 ( .A(\register[3][8] ), .B(n2092), .S0(n936), .Y(n1163) );
  CLKMX2X2 U2081 ( .A(\register[3][9] ), .B(n2097), .S0(n936), .Y(n1162) );
  CLKMX2X2 U2082 ( .A(\register[3][10] ), .B(n2102), .S0(n936), .Y(n1161) );
  CLKMX2X2 U2083 ( .A(\register[3][11] ), .B(n2107), .S0(n936), .Y(n1160) );
  CLKMX2X2 U2084 ( .A(\register[3][12] ), .B(n2112), .S0(n936), .Y(n1159) );
  CLKMX2X2 U2085 ( .A(\register[3][13] ), .B(n2117), .S0(n936), .Y(n1158) );
  CLKMX2X2 U2086 ( .A(\register[3][14] ), .B(n2122), .S0(n936), .Y(n1157) );
  CLKMX2X2 U2087 ( .A(\register[3][15] ), .B(n2127), .S0(n936), .Y(n1156) );
  CLKMX2X2 U2088 ( .A(\register[3][16] ), .B(n2132), .S0(n936), .Y(n1155) );
  CLKMX2X2 U2089 ( .A(\register[3][17] ), .B(n2137), .S0(n936), .Y(n1154) );
  CLKMX2X2 U2090 ( .A(\register[3][18] ), .B(n2142), .S0(n936), .Y(n1153) );
  CLKMX2X2 U2091 ( .A(\register[3][19] ), .B(n2147), .S0(n936), .Y(n1152) );
  CLKMX2X2 U2092 ( .A(\register[3][20] ), .B(n2152), .S0(n935), .Y(n1151) );
  CLKMX2X2 U2093 ( .A(\register[3][21] ), .B(n2157), .S0(n935), .Y(n1150) );
  CLKMX2X2 U2094 ( .A(\register[3][22] ), .B(n2162), .S0(n935), .Y(n1149) );
  CLKMX2X2 U2095 ( .A(\register[3][23] ), .B(n2167), .S0(n935), .Y(n1148) );
  CLKMX2X2 U2096 ( .A(\register[3][24] ), .B(n2172), .S0(n935), .Y(n1147) );
  CLKMX2X2 U2097 ( .A(\register[3][25] ), .B(n2177), .S0(n935), .Y(n1146) );
  CLKMX2X2 U2098 ( .A(\register[3][26] ), .B(n2182), .S0(n935), .Y(n1145) );
  CLKMX2X2 U2099 ( .A(\register[3][27] ), .B(n2187), .S0(n935), .Y(n1144) );
  CLKMX2X2 U2100 ( .A(\register[3][28] ), .B(n2192), .S0(n935), .Y(n1143) );
  CLKMX2X2 U2101 ( .A(\register[3][29] ), .B(n2197), .S0(n935), .Y(n1142) );
  CLKMX2X2 U2102 ( .A(\register[3][30] ), .B(n2202), .S0(n935), .Y(n1141) );
  CLKMX2X2 U2103 ( .A(\register[3][31] ), .B(n2205), .S0(n935), .Y(n1140) );
  CLKMX2X2 U2104 ( .A(\register[2][8] ), .B(n2092), .S0(n933), .Y(n1131) );
  CLKMX2X2 U2105 ( .A(\register[2][9] ), .B(n2097), .S0(n933), .Y(n1130) );
  CLKMX2X2 U2106 ( .A(\register[2][10] ), .B(n2102), .S0(n933), .Y(n1129) );
  CLKMX2X2 U2107 ( .A(\register[2][11] ), .B(n2107), .S0(n933), .Y(n1128) );
  CLKMX2X2 U2108 ( .A(\register[2][12] ), .B(n2112), .S0(n933), .Y(n1127) );
  CLKMX2X2 U2109 ( .A(\register[2][13] ), .B(n2117), .S0(n933), .Y(n1126) );
  CLKMX2X2 U2110 ( .A(\register[2][14] ), .B(n2122), .S0(n933), .Y(n1125) );
  CLKMX2X2 U2111 ( .A(\register[2][15] ), .B(n2127), .S0(n933), .Y(n1124) );
  CLKMX2X2 U2112 ( .A(\register[2][16] ), .B(n2132), .S0(n933), .Y(n1123) );
  CLKMX2X2 U2113 ( .A(\register[2][17] ), .B(n2137), .S0(n933), .Y(n1122) );
  CLKMX2X2 U2114 ( .A(\register[2][18] ), .B(n2142), .S0(n933), .Y(n1121) );
  CLKMX2X2 U2115 ( .A(\register[2][19] ), .B(n2147), .S0(n933), .Y(n1120) );
  CLKMX2X2 U2116 ( .A(\register[2][20] ), .B(n2152), .S0(n932), .Y(n1119) );
  CLKMX2X2 U2117 ( .A(\register[2][21] ), .B(n2157), .S0(n932), .Y(n1118) );
  CLKMX2X2 U2118 ( .A(\register[2][22] ), .B(n2162), .S0(n932), .Y(n1117) );
  CLKMX2X2 U2119 ( .A(\register[2][23] ), .B(n2167), .S0(n932), .Y(n1116) );
  CLKMX2X2 U2120 ( .A(\register[2][24] ), .B(n2172), .S0(n932), .Y(n1115) );
  CLKMX2X2 U2121 ( .A(\register[2][25] ), .B(n2177), .S0(n932), .Y(n1114) );
  CLKMX2X2 U2122 ( .A(\register[2][26] ), .B(n2182), .S0(n932), .Y(n1113) );
  CLKMX2X2 U2123 ( .A(\register[2][27] ), .B(n2187), .S0(n932), .Y(n1112) );
  CLKMX2X2 U2124 ( .A(\register[2][28] ), .B(n2192), .S0(n932), .Y(n1111) );
  CLKMX2X2 U2125 ( .A(\register[2][29] ), .B(n2197), .S0(n932), .Y(n1110) );
  CLKMX2X2 U2126 ( .A(\register[2][30] ), .B(n2202), .S0(n932), .Y(n1109) );
  CLKMX2X2 U2127 ( .A(\register[2][31] ), .B(n2205), .S0(n932), .Y(n1108) );
  CLKMX2X2 U2128 ( .A(\register[1][8] ), .B(n2092), .S0(n930), .Y(n1099) );
  CLKMX2X2 U2129 ( .A(\register[1][9] ), .B(n2097), .S0(n930), .Y(n1098) );
  CLKMX2X2 U2130 ( .A(\register[1][10] ), .B(n2102), .S0(n930), .Y(n1097) );
  CLKMX2X2 U2131 ( .A(\register[1][11] ), .B(n2107), .S0(n930), .Y(n1096) );
  CLKMX2X2 U2132 ( .A(\register[1][12] ), .B(n2112), .S0(n930), .Y(n1095) );
  CLKMX2X2 U2133 ( .A(\register[1][13] ), .B(n2117), .S0(n930), .Y(n1094) );
  CLKMX2X2 U2134 ( .A(\register[1][14] ), .B(n2122), .S0(n930), .Y(n1093) );
  CLKMX2X2 U2135 ( .A(\register[1][15] ), .B(n2127), .S0(n930), .Y(n1092) );
  CLKMX2X2 U2136 ( .A(\register[1][16] ), .B(n2132), .S0(n930), .Y(n1091) );
  CLKMX2X2 U2137 ( .A(\register[1][17] ), .B(n2137), .S0(n930), .Y(n1090) );
  CLKMX2X2 U2138 ( .A(\register[1][18] ), .B(n2142), .S0(n930), .Y(n1089) );
  CLKMX2X2 U2139 ( .A(\register[1][19] ), .B(n2147), .S0(n930), .Y(n1088) );
  CLKMX2X2 U2140 ( .A(\register[1][20] ), .B(n2152), .S0(n929), .Y(n1087) );
  CLKMX2X2 U2141 ( .A(\register[1][21] ), .B(n2157), .S0(n929), .Y(n1086) );
  CLKMX2X2 U2142 ( .A(\register[1][22] ), .B(n2162), .S0(n929), .Y(n1085) );
  CLKMX2X2 U2143 ( .A(\register[1][23] ), .B(n2167), .S0(n929), .Y(n1084) );
  CLKMX2X2 U2144 ( .A(\register[1][24] ), .B(n2172), .S0(n929), .Y(n1083) );
  CLKMX2X2 U2145 ( .A(\register[1][25] ), .B(n2177), .S0(n929), .Y(n1082) );
  CLKMX2X2 U2146 ( .A(\register[1][26] ), .B(n2182), .S0(n929), .Y(n1081) );
  CLKMX2X2 U2147 ( .A(\register[1][27] ), .B(n2187), .S0(n929), .Y(n1080) );
  CLKMX2X2 U2148 ( .A(\register[1][28] ), .B(n2192), .S0(n929), .Y(n1079) );
  CLKMX2X2 U2149 ( .A(\register[1][29] ), .B(n2197), .S0(n929), .Y(n1078) );
  CLKMX2X2 U2150 ( .A(\register[1][30] ), .B(n2202), .S0(n929), .Y(n1077) );
  CLKMX2X2 U2151 ( .A(\register[1][31] ), .B(n2205), .S0(n929), .Y(n1076) );
  CLKMX2X2 U2152 ( .A(\register[0][8] ), .B(n2092), .S0(n927), .Y(n1067) );
  CLKMX2X2 U2153 ( .A(\register[0][9] ), .B(n2097), .S0(n927), .Y(n1066) );
  CLKMX2X2 U2154 ( .A(\register[0][10] ), .B(n2102), .S0(n927), .Y(n1065) );
  CLKMX2X2 U2155 ( .A(\register[0][11] ), .B(n2107), .S0(n927), .Y(n1064) );
  CLKMX2X2 U2156 ( .A(\register[0][12] ), .B(n2112), .S0(n927), .Y(n1063) );
  CLKMX2X2 U2157 ( .A(\register[0][13] ), .B(n2117), .S0(n927), .Y(n1062) );
  CLKMX2X2 U2158 ( .A(\register[0][14] ), .B(n2122), .S0(n927), .Y(n1061) );
  CLKMX2X2 U2159 ( .A(\register[0][15] ), .B(n2127), .S0(n927), .Y(n1060) );
  CLKMX2X2 U2160 ( .A(\register[0][16] ), .B(n2132), .S0(n927), .Y(n1059) );
  CLKMX2X2 U2161 ( .A(\register[0][17] ), .B(n2137), .S0(n927), .Y(n1058) );
  CLKMX2X2 U2162 ( .A(\register[0][18] ), .B(n2142), .S0(n927), .Y(n1057) );
  CLKMX2X2 U2163 ( .A(\register[0][19] ), .B(n2147), .S0(n927), .Y(n1056) );
  CLKMX2X2 U2164 ( .A(\register[0][20] ), .B(n2152), .S0(n926), .Y(n1055) );
  CLKMX2X2 U2165 ( .A(\register[0][21] ), .B(n2157), .S0(n926), .Y(n1054) );
  CLKMX2X2 U2166 ( .A(\register[0][22] ), .B(n2162), .S0(n926), .Y(n1053) );
  CLKMX2X2 U2167 ( .A(\register[0][23] ), .B(n2167), .S0(n926), .Y(n1052) );
  CLKMX2X2 U2168 ( .A(\register[0][24] ), .B(n2172), .S0(n926), .Y(n1051) );
  CLKMX2X2 U2169 ( .A(\register[0][25] ), .B(n2177), .S0(n926), .Y(n1050) );
  CLKMX2X2 U2170 ( .A(\register[0][26] ), .B(n2182), .S0(n926), .Y(n1049) );
  CLKMX2X2 U2171 ( .A(\register[0][27] ), .B(n2187), .S0(n926), .Y(n1048) );
  CLKMX2X2 U2172 ( .A(\register[0][28] ), .B(n2192), .S0(n926), .Y(n1047) );
  CLKMX2X2 U2173 ( .A(\register[0][29] ), .B(n2197), .S0(n926), .Y(n1046) );
  CLKMX2X2 U2174 ( .A(\register[0][30] ), .B(n2202), .S0(n926), .Y(n1045) );
  CLKMX2X2 U2175 ( .A(\register[0][31] ), .B(n2205), .S0(n926), .Y(n1044) );
  CLKMX2X2 U2176 ( .A(n66), .B(n67), .S0(n395), .Y(ReadData1_o[14]) );
  MXI4X1 U2177 ( .A(n254), .B(n252), .C(n253), .D(n251), .S0(n402), .S1(n410), 
        .Y(n66) );
  MXI4X1 U2178 ( .A(n250), .B(n248), .C(n249), .D(n247), .S0(n402), .S1(n410), 
        .Y(n67) );
  CLKMX2X2 U2179 ( .A(n68), .B(n71), .S0(n395), .Y(ReadData1_o[17]) );
  MXI4X1 U2180 ( .A(n279), .B(n277), .C(n278), .D(n276), .S0(n402), .S1(n410), 
        .Y(n68) );
  MXI4X1 U2181 ( .A(n275), .B(n272), .C(n273), .D(n271), .S0(n402), .S1(n410), 
        .Y(n71) );
  CLKMX2X2 U2182 ( .A(n72), .B(n73), .S0(n395), .Y(ReadData1_o[16]) );
  MXI4X1 U2183 ( .A(n270), .B(n268), .C(n269), .D(n267), .S0(n402), .S1(n410), 
        .Y(n72) );
  MXI4X1 U2184 ( .A(n266), .B(n264), .C(n265), .D(n263), .S0(n402), .S1(n410), 
        .Y(n73) );
  MX4X1 U2185 ( .A(n295), .B(n293), .C(n294), .D(n292), .S0(n402), .S1(n411), 
        .Y(n111) );
  MX4X1 U2186 ( .A(n291), .B(n289), .C(n290), .D(n288), .S0(n402), .S1(n411), 
        .Y(n112) );
  MXI4X1 U2187 ( .A(\register[0][19] ), .B(\register[1][19] ), .C(
        \register[2][19] ), .D(\register[3][19] ), .S0(n487), .S1(n446), .Y(
        n295) );
  MX4X1 U2188 ( .A(n229), .B(n227), .C(n228), .D(n226), .S0(n401), .S1(n409), 
        .Y(n100) );
  MX4X1 U2189 ( .A(n225), .B(n223), .C(n224), .D(n222), .S0(n401), .S1(n409), 
        .Y(n101) );
  MXI4X1 U2190 ( .A(\register[0][11] ), .B(\register[1][11] ), .C(
        \register[2][11] ), .D(\register[3][11] ), .S0(n482), .S1(n441), .Y(
        n229) );
  MX4X1 U2191 ( .A(n246), .B(n244), .C(n245), .D(n243), .S0(n401), .S1(n410), 
        .Y(n105) );
  MX4X1 U2192 ( .A(n242), .B(n239), .C(n241), .D(n238), .S0(n401), .S1(n410), 
        .Y(n106) );
  MXI4X1 U2193 ( .A(\register[0][13] ), .B(\register[1][13] ), .C(
        \register[2][13] ), .D(\register[3][13] ), .S0(n483), .S1(n442), .Y(
        n246) );
  MX4X1 U2194 ( .A(n312), .B(n310), .C(n311), .D(n309), .S0(n403), .S1(n411), 
        .Y(n115) );
  MX4X1 U2195 ( .A(n307), .B(n305), .C(n306), .D(n304), .S0(n403), .S1(n411), 
        .Y(n116) );
  MXI4X1 U2196 ( .A(\register[8][21] ), .B(\register[9][21] ), .C(
        \register[10][21] ), .D(\register[11][21] ), .S0(n489), .S1(n448), .Y(
        n310) );
  MX4X1 U2197 ( .A(n221), .B(n219), .C(n220), .D(n218), .S0(n401), .S1(n409), 
        .Y(n98) );
  MX4X1 U2198 ( .A(n217), .B(n215), .C(n216), .D(n214), .S0(n401), .S1(n409), 
        .Y(n99) );
  MXI4X1 U2199 ( .A(\register[0][10] ), .B(\register[1][10] ), .C(
        \register[2][10] ), .D(\register[3][10] ), .S0(n481), .S1(n440), .Y(
        n221) );
  MX4X1 U2200 ( .A(n237), .B(n235), .C(n236), .D(n234), .S0(n401), .S1(n410), 
        .Y(n102) );
  MX4X1 U2201 ( .A(n233), .B(n231), .C(n232), .D(n230), .S0(n401), .S1(n409), 
        .Y(n103) );
  MXI4X1 U2202 ( .A(\register[0][12] ), .B(\register[1][12] ), .C(
        \register[2][12] ), .D(\register[3][12] ), .S0(n483), .S1(n442), .Y(
        n237) );
  MX4X1 U2203 ( .A(n303), .B(n301), .C(n302), .D(n300), .S0(n403), .S1(n411), 
        .Y(n113) );
  MX4X1 U2204 ( .A(n299), .B(n297), .C(n298), .D(n296), .S0(n403), .S1(n411), 
        .Y(n114) );
  MXI4X1 U2205 ( .A(\register[0][20] ), .B(\register[1][20] ), .C(
        \register[2][20] ), .D(\register[3][20] ), .S0(n488), .S1(n447), .Y(
        n303) );
  MX4X1 U2206 ( .A(n262), .B(n260), .C(n261), .D(n259), .S0(n402), .S1(n410), 
        .Y(n107) );
  MX4X1 U2207 ( .A(n258), .B(n256), .C(n257), .D(n255), .S0(n402), .S1(n410), 
        .Y(n108) );
  MXI4X1 U2208 ( .A(\register[0][15] ), .B(\register[1][15] ), .C(
        \register[2][15] ), .D(\register[3][15] ), .S0(n485), .S1(n444), .Y(
        n262) );
  MX4X1 U2209 ( .A(n213), .B(n211), .C(n212), .D(n210), .S0(n401), .S1(n409), 
        .Y(n96) );
  MX4X1 U2210 ( .A(n209), .B(n207), .C(n208), .D(n205), .S0(n401), .S1(n409), 
        .Y(n97) );
  MXI4X1 U2211 ( .A(\register[0][9] ), .B(\register[1][9] ), .C(
        \register[2][9] ), .D(\register[3][9] ), .S0(n481), .S1(n440), .Y(n213) );
  MX4X1 U2212 ( .A(n287), .B(n285), .C(n286), .D(n284), .S0(n402), .S1(n410), 
        .Y(n109) );
  MX4X1 U2213 ( .A(n283), .B(n281), .C(n282), .D(n280), .S0(n402), .S1(n410), 
        .Y(n110) );
  MXI4X1 U2214 ( .A(\register[0][18] ), .B(\register[1][18] ), .C(
        \register[2][18] ), .D(\register[3][18] ), .S0(n487), .S1(n446), .Y(
        n287) );
  MXI4X1 U2215 ( .A(\register[20][9] ), .B(\register[21][9] ), .C(
        \register[22][9] ), .D(\register[23][9] ), .S0(n480), .S1(n439), .Y(
        n208) );
  MXI4X1 U2216 ( .A(\register[4][9] ), .B(\register[5][9] ), .C(
        \register[6][9] ), .D(\register[7][9] ), .S0(n481), .S1(n440), .Y(n212) );
  MXI4X1 U2217 ( .A(\register[20][11] ), .B(\register[21][11] ), .C(
        \register[22][11] ), .D(\register[23][11] ), .S0(n482), .S1(n441), .Y(
        n224) );
  MXI4X1 U2218 ( .A(\register[4][11] ), .B(\register[5][11] ), .C(
        \register[6][11] ), .D(\register[7][11] ), .S0(n482), .S1(n441), .Y(
        n228) );
  MXI4X1 U2219 ( .A(\register[20][13] ), .B(\register[21][13] ), .C(
        \register[22][13] ), .D(\register[23][13] ), .S0(n483), .S1(n442), .Y(
        n241) );
  MXI4X1 U2220 ( .A(\register[4][13] ), .B(\register[5][13] ), .C(
        \register[6][13] ), .D(\register[7][13] ), .S0(n483), .S1(n442), .Y(
        n245) );
  MXI4X1 U2221 ( .A(\register[20][15] ), .B(\register[21][15] ), .C(
        \register[22][15] ), .D(\register[23][15] ), .S0(n484), .S1(n443), .Y(
        n257) );
  MXI4X1 U2222 ( .A(\register[4][15] ), .B(\register[5][15] ), .C(
        \register[6][15] ), .D(\register[7][15] ), .S0(n485), .S1(n444), .Y(
        n261) );
  MXI4X1 U2223 ( .A(\register[20][17] ), .B(\register[21][17] ), .C(
        \register[22][17] ), .D(\register[23][17] ), .S0(n486), .S1(n445), .Y(
        n273) );
  MXI4X1 U2224 ( .A(\register[4][17] ), .B(\register[5][17] ), .C(
        \register[6][17] ), .D(\register[7][17] ), .S0(n486), .S1(n445), .Y(
        n278) );
  MXI4X1 U2225 ( .A(\register[20][19] ), .B(\register[21][19] ), .C(
        \register[22][19] ), .D(\register[23][19] ), .S0(n487), .S1(n446), .Y(
        n290) );
  MXI4X1 U2226 ( .A(\register[4][19] ), .B(\register[5][19] ), .C(
        \register[6][19] ), .D(\register[7][19] ), .S0(n487), .S1(n446), .Y(
        n294) );
  MXI4X1 U2227 ( .A(\register[20][21] ), .B(\register[21][21] ), .C(
        \register[22][21] ), .D(\register[23][21] ), .S0(n488), .S1(n447), .Y(
        n306) );
  MXI4X1 U2228 ( .A(\register[4][21] ), .B(\register[5][21] ), .C(
        \register[6][21] ), .D(\register[7][21] ), .S0(n489), .S1(n448), .Y(
        n311) );
  MXI4X1 U2229 ( .A(\register[20][10] ), .B(\register[21][10] ), .C(
        \register[22][10] ), .D(\register[23][10] ), .S0(n481), .S1(n440), .Y(
        n216) );
  MXI4X1 U2230 ( .A(\register[4][10] ), .B(\register[5][10] ), .C(
        \register[6][10] ), .D(\register[7][10] ), .S0(n481), .S1(n440), .Y(
        n220) );
  MXI4X1 U2231 ( .A(\register[20][12] ), .B(\register[21][12] ), .C(
        \register[22][12] ), .D(\register[23][12] ), .S0(n482), .S1(n441), .Y(
        n232) );
  MXI4X1 U2232 ( .A(\register[4][12] ), .B(\register[5][12] ), .C(
        \register[6][12] ), .D(\register[7][12] ), .S0(n483), .S1(n442), .Y(
        n236) );
  MXI4X1 U2233 ( .A(\register[20][14] ), .B(\register[21][14] ), .C(
        \register[22][14] ), .D(\register[23][14] ), .S0(n484), .S1(n443), .Y(
        n249) );
  MXI4X1 U2234 ( .A(\register[4][14] ), .B(\register[5][14] ), .C(
        \register[6][14] ), .D(\register[7][14] ), .S0(n484), .S1(n443), .Y(
        n253) );
  MXI4X1 U2235 ( .A(\register[20][16] ), .B(\register[21][16] ), .C(
        \register[22][16] ), .D(\register[23][16] ), .S0(n485), .S1(n444), .Y(
        n265) );
  MXI4X1 U2236 ( .A(\register[4][16] ), .B(\register[5][16] ), .C(
        \register[6][16] ), .D(\register[7][16] ), .S0(n485), .S1(n444), .Y(
        n269) );
  MXI4X1 U2237 ( .A(\register[20][18] ), .B(\register[21][18] ), .C(
        \register[22][18] ), .D(\register[23][18] ), .S0(n486), .S1(n445), .Y(
        n282) );
  MXI4X1 U2238 ( .A(\register[4][18] ), .B(\register[5][18] ), .C(
        \register[6][18] ), .D(\register[7][18] ), .S0(n487), .S1(n446), .Y(
        n286) );
  MXI4X1 U2239 ( .A(\register[20][20] ), .B(\register[21][20] ), .C(
        \register[22][20] ), .D(\register[23][20] ), .S0(n488), .S1(n447), .Y(
        n298) );
  MXI4X1 U2240 ( .A(\register[4][20] ), .B(\register[5][20] ), .C(
        \register[6][20] ), .D(\register[7][20] ), .S0(n488), .S1(n447), .Y(
        n302) );
  MXI4X1 U2241 ( .A(\register[16][9] ), .B(\register[17][9] ), .C(
        \register[18][9] ), .D(\register[19][9] ), .S0(n480), .S1(n439), .Y(
        n209) );
  MXI4X1 U2242 ( .A(\register[16][11] ), .B(\register[17][11] ), .C(
        \register[18][11] ), .D(\register[19][11] ), .S0(n482), .S1(n441), .Y(
        n225) );
  MXI4X1 U2243 ( .A(\register[16][13] ), .B(\register[17][13] ), .C(
        \register[18][13] ), .D(\register[19][13] ), .S0(n483), .S1(n442), .Y(
        n242) );
  MXI4X1 U2244 ( .A(\register[16][15] ), .B(\register[17][15] ), .C(
        \register[18][15] ), .D(\register[19][15] ), .S0(n484), .S1(n443), .Y(
        n258) );
  MXI4X1 U2245 ( .A(\register[16][17] ), .B(\register[17][17] ), .C(
        \register[18][17] ), .D(\register[19][17] ), .S0(n486), .S1(n445), .Y(
        n275) );
  MXI4X1 U2246 ( .A(\register[16][19] ), .B(\register[17][19] ), .C(
        \register[18][19] ), .D(\register[19][19] ), .S0(n487), .S1(n446), .Y(
        n291) );
  MXI4X1 U2247 ( .A(\register[16][21] ), .B(\register[17][21] ), .C(
        \register[18][21] ), .D(\register[19][21] ), .S0(n488), .S1(n447), .Y(
        n307) );
  MXI4X1 U2248 ( .A(\register[0][21] ), .B(\register[1][21] ), .C(
        \register[2][21] ), .D(\register[3][21] ), .S0(n489), .S1(n448), .Y(
        n312) );
  MXI4X1 U2249 ( .A(\register[16][10] ), .B(\register[17][10] ), .C(
        \register[18][10] ), .D(\register[19][10] ), .S0(n481), .S1(n440), .Y(
        n217) );
  MXI4X1 U2250 ( .A(\register[16][12] ), .B(\register[17][12] ), .C(
        \register[18][12] ), .D(\register[19][12] ), .S0(n482), .S1(n441), .Y(
        n233) );
  MXI4X1 U2251 ( .A(\register[16][14] ), .B(\register[17][14] ), .C(
        \register[18][14] ), .D(\register[19][14] ), .S0(n484), .S1(n443), .Y(
        n250) );
  MXI4X1 U2252 ( .A(\register[16][16] ), .B(\register[17][16] ), .C(
        \register[18][16] ), .D(\register[19][16] ), .S0(n485), .S1(n444), .Y(
        n266) );
  MXI4X1 U2253 ( .A(\register[16][18] ), .B(\register[17][18] ), .C(
        \register[18][18] ), .D(\register[19][18] ), .S0(n486), .S1(n445), .Y(
        n283) );
  MXI4X1 U2254 ( .A(\register[16][20] ), .B(\register[17][20] ), .C(
        \register[18][20] ), .D(\register[19][20] ), .S0(n488), .S1(n447), .Y(
        n299) );
  MXI4X1 U2255 ( .A(\register[28][9] ), .B(\register[29][9] ), .C(
        \register[30][9] ), .D(\register[31][9] ), .S0(n480), .S1(n439), .Y(
        n205) );
  MXI4X1 U2256 ( .A(\register[12][9] ), .B(\register[13][9] ), .C(
        \register[14][9] ), .D(\register[15][9] ), .S0(n481), .S1(n440), .Y(
        n210) );
  MXI4X1 U2257 ( .A(\register[28][11] ), .B(\register[29][11] ), .C(
        \register[30][11] ), .D(\register[31][11] ), .S0(n482), .S1(n441), .Y(
        n222) );
  MXI4X1 U2258 ( .A(\register[12][11] ), .B(\register[13][11] ), .C(
        \register[14][11] ), .D(\register[15][11] ), .S0(n482), .S1(n441), .Y(
        n226) );
  MXI4X1 U2259 ( .A(\register[28][13] ), .B(\register[29][13] ), .C(
        \register[30][13] ), .D(\register[31][13] ), .S0(n483), .S1(n442), .Y(
        n238) );
  MXI4X1 U2260 ( .A(\register[12][13] ), .B(\register[13][13] ), .C(
        \register[14][13] ), .D(\register[15][13] ), .S0(n483), .S1(n442), .Y(
        n243) );
  MXI4X1 U2261 ( .A(\register[28][15] ), .B(\register[29][15] ), .C(
        \register[30][15] ), .D(\register[31][15] ), .S0(n484), .S1(n443), .Y(
        n255) );
  MXI4X1 U2262 ( .A(\register[12][15] ), .B(\register[13][15] ), .C(
        \register[14][15] ), .D(\register[15][15] ), .S0(n485), .S1(n444), .Y(
        n259) );
  MXI4X1 U2263 ( .A(\register[28][17] ), .B(\register[29][17] ), .C(
        \register[30][17] ), .D(\register[31][17] ), .S0(n486), .S1(n445), .Y(
        n271) );
  MXI4X1 U2264 ( .A(\register[12][17] ), .B(\register[13][17] ), .C(
        \register[14][17] ), .D(\register[15][17] ), .S0(n486), .S1(n445), .Y(
        n276) );
  MXI4X1 U2265 ( .A(\register[28][19] ), .B(\register[29][19] ), .C(
        \register[30][19] ), .D(\register[31][19] ), .S0(n487), .S1(n446), .Y(
        n288) );
  MXI4X1 U2266 ( .A(\register[12][19] ), .B(\register[13][19] ), .C(
        \register[14][19] ), .D(\register[15][19] ), .S0(n487), .S1(n446), .Y(
        n292) );
  MXI4X1 U2267 ( .A(\register[28][21] ), .B(\register[29][21] ), .C(
        \register[30][21] ), .D(\register[31][21] ), .S0(n488), .S1(n447), .Y(
        n304) );
  MXI4X1 U2268 ( .A(\register[12][21] ), .B(\register[13][21] ), .C(
        \register[14][21] ), .D(\register[15][21] ), .S0(n489), .S1(n448), .Y(
        n309) );
  MXI4X1 U2269 ( .A(\register[28][10] ), .B(\register[29][10] ), .C(
        \register[30][10] ), .D(\register[31][10] ), .S0(n481), .S1(n440), .Y(
        n214) );
  MXI4X1 U2270 ( .A(\register[12][10] ), .B(\register[13][10] ), .C(
        \register[14][10] ), .D(\register[15][10] ), .S0(n481), .S1(n440), .Y(
        n218) );
  MXI4X1 U2271 ( .A(\register[28][12] ), .B(\register[29][12] ), .C(
        \register[30][12] ), .D(\register[31][12] ), .S0(n482), .S1(n441), .Y(
        n230) );
  MXI4X1 U2272 ( .A(\register[12][12] ), .B(\register[13][12] ), .C(
        \register[14][12] ), .D(\register[15][12] ), .S0(n483), .S1(n442), .Y(
        n234) );
  MXI4X1 U2273 ( .A(\register[28][14] ), .B(\register[29][14] ), .C(
        \register[30][14] ), .D(\register[31][14] ), .S0(n484), .S1(n443), .Y(
        n247) );
  MXI4X1 U2274 ( .A(\register[12][14] ), .B(\register[13][14] ), .C(
        \register[14][14] ), .D(\register[15][14] ), .S0(n484), .S1(n443), .Y(
        n251) );
  MXI4X1 U2275 ( .A(\register[28][16] ), .B(\register[29][16] ), .C(
        \register[30][16] ), .D(\register[31][16] ), .S0(n485), .S1(n444), .Y(
        n263) );
  MXI4X1 U2276 ( .A(\register[12][16] ), .B(\register[13][16] ), .C(
        \register[14][16] ), .D(\register[15][16] ), .S0(n485), .S1(n444), .Y(
        n267) );
  MXI4X1 U2277 ( .A(\register[28][18] ), .B(\register[29][18] ), .C(
        \register[30][18] ), .D(\register[31][18] ), .S0(n486), .S1(n445), .Y(
        n280) );
  MXI4X1 U2278 ( .A(\register[12][18] ), .B(\register[13][18] ), .C(
        \register[14][18] ), .D(\register[15][18] ), .S0(n487), .S1(n446), .Y(
        n284) );
  MXI4X1 U2279 ( .A(\register[28][20] ), .B(\register[29][20] ), .C(
        \register[30][20] ), .D(\register[31][20] ), .S0(n488), .S1(n447), .Y(
        n296) );
  MXI4X1 U2280 ( .A(\register[12][20] ), .B(\register[13][20] ), .C(
        \register[14][20] ), .D(\register[15][20] ), .S0(n488), .S1(n447), .Y(
        n300) );
  MXI4X1 U2281 ( .A(\register[24][9] ), .B(\register[25][9] ), .C(
        \register[26][9] ), .D(\register[27][9] ), .S0(n480), .S1(n439), .Y(
        n207) );
  MXI4X1 U2282 ( .A(\register[8][9] ), .B(\register[9][9] ), .C(
        \register[10][9] ), .D(\register[11][9] ), .S0(n481), .S1(n440), .Y(
        n211) );
  MXI4X1 U2283 ( .A(\register[24][11] ), .B(\register[25][11] ), .C(
        \register[26][11] ), .D(\register[27][11] ), .S0(n482), .S1(n441), .Y(
        n223) );
  MXI4X1 U2284 ( .A(\register[8][11] ), .B(\register[9][11] ), .C(
        \register[10][11] ), .D(\register[11][11] ), .S0(n482), .S1(n441), .Y(
        n227) );
  MXI4X1 U2285 ( .A(\register[24][13] ), .B(\register[25][13] ), .C(
        \register[26][13] ), .D(\register[27][13] ), .S0(n483), .S1(n442), .Y(
        n239) );
  MXI4X1 U2286 ( .A(\register[8][13] ), .B(\register[9][13] ), .C(
        \register[10][13] ), .D(\register[11][13] ), .S0(n483), .S1(n442), .Y(
        n244) );
  MXI4X1 U2287 ( .A(\register[24][15] ), .B(\register[25][15] ), .C(
        \register[26][15] ), .D(\register[27][15] ), .S0(n484), .S1(n443), .Y(
        n256) );
  MXI4X1 U2288 ( .A(\register[8][15] ), .B(\register[9][15] ), .C(
        \register[10][15] ), .D(\register[11][15] ), .S0(n485), .S1(n444), .Y(
        n260) );
  MXI4X1 U2289 ( .A(\register[24][17] ), .B(\register[25][17] ), .C(
        \register[26][17] ), .D(\register[27][17] ), .S0(n486), .S1(n445), .Y(
        n272) );
  MXI4X1 U2290 ( .A(\register[8][17] ), .B(\register[9][17] ), .C(
        \register[10][17] ), .D(\register[11][17] ), .S0(n486), .S1(n445), .Y(
        n277) );
  MXI4X1 U2291 ( .A(\register[24][19] ), .B(\register[25][19] ), .C(
        \register[26][19] ), .D(\register[27][19] ), .S0(n487), .S1(n446), .Y(
        n289) );
  MXI4X1 U2292 ( .A(\register[8][19] ), .B(\register[9][19] ), .C(
        \register[10][19] ), .D(\register[11][19] ), .S0(n487), .S1(n446), .Y(
        n293) );
  MXI4X1 U2293 ( .A(\register[24][21] ), .B(\register[25][21] ), .C(
        \register[26][21] ), .D(\register[27][21] ), .S0(n488), .S1(n447), .Y(
        n305) );
  MXI4X1 U2294 ( .A(\register[24][10] ), .B(\register[25][10] ), .C(
        \register[26][10] ), .D(\register[27][10] ), .S0(n481), .S1(n440), .Y(
        n215) );
  MXI4X1 U2295 ( .A(\register[8][10] ), .B(\register[9][10] ), .C(
        \register[10][10] ), .D(\register[11][10] ), .S0(n481), .S1(n440), .Y(
        n219) );
  MXI4X1 U2296 ( .A(\register[24][12] ), .B(\register[25][12] ), .C(
        \register[26][12] ), .D(\register[27][12] ), .S0(n482), .S1(n441), .Y(
        n231) );
  MXI4X1 U2297 ( .A(\register[8][12] ), .B(\register[9][12] ), .C(
        \register[10][12] ), .D(\register[11][12] ), .S0(n483), .S1(n442), .Y(
        n235) );
  MXI4X1 U2298 ( .A(\register[24][14] ), .B(\register[25][14] ), .C(
        \register[26][14] ), .D(\register[27][14] ), .S0(n484), .S1(n443), .Y(
        n248) );
  MXI4X1 U2299 ( .A(\register[8][14] ), .B(\register[9][14] ), .C(
        \register[10][14] ), .D(\register[11][14] ), .S0(n484), .S1(n443), .Y(
        n252) );
  MXI4X1 U2300 ( .A(\register[24][16] ), .B(\register[25][16] ), .C(
        \register[26][16] ), .D(\register[27][16] ), .S0(n485), .S1(n444), .Y(
        n264) );
  MXI4X1 U2301 ( .A(\register[8][16] ), .B(\register[9][16] ), .C(
        \register[10][16] ), .D(\register[11][16] ), .S0(n485), .S1(n444), .Y(
        n268) );
  MXI4X1 U2302 ( .A(\register[24][18] ), .B(\register[25][18] ), .C(
        \register[26][18] ), .D(\register[27][18] ), .S0(n486), .S1(n445), .Y(
        n281) );
  MXI4X1 U2303 ( .A(\register[8][18] ), .B(\register[9][18] ), .C(
        \register[10][18] ), .D(\register[11][18] ), .S0(n487), .S1(n446), .Y(
        n285) );
  MXI4X1 U2304 ( .A(\register[24][20] ), .B(\register[25][20] ), .C(
        \register[26][20] ), .D(\register[27][20] ), .S0(n488), .S1(n447), .Y(
        n297) );
  MXI4X1 U2305 ( .A(\register[8][20] ), .B(\register[9][20] ), .C(
        \register[10][20] ), .D(\register[11][20] ), .S0(n488), .S1(n447), .Y(
        n301) );
  CLKMX2X2 U2306 ( .A(n74), .B(n75), .S0(n396), .Y(ReadData1_o[22]) );
  MXI4X1 U2307 ( .A(n320), .B(n318), .C(n319), .D(n317), .S0(n403), .S1(n411), 
        .Y(n74) );
  MXI4X1 U2308 ( .A(n316), .B(n314), .C(n315), .D(n313), .S0(n403), .S1(n411), 
        .Y(n75) );
  MX4X1 U2309 ( .A(n373), .B(n371), .C(n372), .D(n370), .S0(n404), .S1(n412), 
        .Y(n126) );
  MX4X1 U2310 ( .A(n377), .B(n375), .C(n376), .D(n374), .S0(n404), .S1(n412), 
        .Y(n125) );
  MXI4X1 U2311 ( .A(\register[28][29] ), .B(\register[29][29] ), .C(
        \register[30][29] ), .D(\register[31][29] ), .S0(n494), .S1(n453), .Y(
        n370) );
  MXI2X1 U2312 ( .A(n129), .B(n130), .S0(n396), .Y(ReadData1_o[31]) );
  MX4X1 U2313 ( .A(n393), .B(n391), .C(n392), .D(n390), .S0(n404), .S1(n412), 
        .Y(n129) );
  MX4X1 U2314 ( .A(n389), .B(n387), .C(n388), .D(n386), .S0(n404), .S1(n412), 
        .Y(n130) );
  MXI4X1 U2315 ( .A(\register[0][31] ), .B(\register[1][31] ), .C(
        \register[2][31] ), .D(\register[3][31] ), .S0(n495), .S1(n454), .Y(
        n393) );
  MXI2X1 U2316 ( .A(n127), .B(n128), .S0(n396), .Y(ReadData1_o[30]) );
  MX4X1 U2317 ( .A(n385), .B(n383), .C(n384), .D(n382), .S0(n404), .S1(n412), 
        .Y(n127) );
  MX4X1 U2318 ( .A(n381), .B(n379), .C(n380), .D(n378), .S0(n404), .S1(n412), 
        .Y(n128) );
  MXI4X1 U2319 ( .A(\register[0][30] ), .B(\register[1][30] ), .C(
        \register[2][30] ), .D(\register[3][30] ), .S0(n495), .S1(n454), .Y(
        n385) );
  MX4X1 U2320 ( .A(n324), .B(n322), .C(n323), .D(n321), .S0(n403), .S1(n411), 
        .Y(n118) );
  MX4X1 U2321 ( .A(n328), .B(n326), .C(n327), .D(n325), .S0(n403), .S1(n411), 
        .Y(n117) );
  MXI4X1 U2322 ( .A(\register[16][23] ), .B(\register[17][23] ), .C(
        \register[18][23] ), .D(\register[19][23] ), .S0(n490), .S1(n449), .Y(
        n324) );
  MX4X1 U2323 ( .A(n357), .B(n355), .C(n356), .D(n354), .S0(n404), .S1(n412), 
        .Y(n122) );
  MX4X1 U2324 ( .A(n361), .B(n359), .C(n360), .D(n358), .S0(n404), .S1(n412), 
        .Y(n121) );
  MXI4X1 U2325 ( .A(\register[28][27] ), .B(\register[29][27] ), .C(
        \register[30][27] ), .D(\register[31][27] ), .S0(n492), .S1(n451), .Y(
        n354) );
  MX4X1 U2326 ( .A(n349), .B(n347), .C(n348), .D(n346), .S0(n404), .S1(n412), 
        .Y(n120) );
  MX4X1 U2327 ( .A(n353), .B(n351), .C(n352), .D(n350), .S0(n404), .S1(n412), 
        .Y(n119) );
  MXI4X1 U2328 ( .A(\register[28][26] ), .B(\register[29][26] ), .C(
        \register[30][26] ), .D(\register[31][26] ), .S0(n492), .S1(n451), .Y(
        n346) );
  MX4X1 U2329 ( .A(n365), .B(n363), .C(n364), .D(n362), .S0(n404), .S1(n412), 
        .Y(n124) );
  MX4X1 U2330 ( .A(n369), .B(n367), .C(n368), .D(n366), .S0(n404), .S1(n412), 
        .Y(n123) );
  MXI4X1 U2331 ( .A(\register[28][28] ), .B(\register[29][28] ), .C(
        \register[30][28] ), .D(\register[31][28] ), .S0(n493), .S1(n452), .Y(
        n362) );
  CLKMX2X2 U2332 ( .A(n76), .B(n77), .S0(n396), .Y(ReadData1_o[25]) );
  MXI4X1 U2333 ( .A(n345), .B(n343), .C(n344), .D(n341), .S0(n403), .S1(n412), 
        .Y(n76) );
  MXI4X1 U2334 ( .A(n340), .B(n338), .C(n339), .D(n337), .S0(n403), .S1(n411), 
        .Y(n77) );
  CLKMX2X2 U2335 ( .A(n78), .B(n79), .S0(n396), .Y(ReadData1_o[24]) );
  MXI4X1 U2336 ( .A(n336), .B(n334), .C(n335), .D(n333), .S0(n403), .S1(n411), 
        .Y(n78) );
  MXI4X1 U2337 ( .A(n332), .B(n330), .C(n331), .D(n329), .S0(n403), .S1(n411), 
        .Y(n79) );
  MXI4X1 U2338 ( .A(\register[4][23] ), .B(\register[5][23] ), .C(
        \register[6][23] ), .D(\register[7][23] ), .S0(n490), .S1(n449), .Y(
        n327) );
  MXI4X1 U2339 ( .A(\register[20][23] ), .B(\register[21][23] ), .C(
        \register[22][23] ), .D(\register[23][23] ), .S0(n490), .S1(n449), .Y(
        n323) );
  MXI4X1 U2340 ( .A(\register[20][25] ), .B(\register[21][25] ), .C(
        \register[22][25] ), .D(\register[23][25] ), .S0(n491), .S1(n450), .Y(
        n339) );
  MXI4X1 U2341 ( .A(\register[4][25] ), .B(\register[5][25] ), .C(
        \register[6][25] ), .D(\register[7][25] ), .S0(n491), .S1(n450), .Y(
        n344) );
  MXI4X1 U2342 ( .A(\register[4][27] ), .B(\register[5][27] ), .C(
        \register[6][27] ), .D(\register[7][27] ), .S0(n493), .S1(n452), .Y(
        n360) );
  MXI4X1 U2343 ( .A(\register[20][27] ), .B(\register[21][27] ), .C(
        \register[22][27] ), .D(\register[23][27] ), .S0(n492), .S1(n451), .Y(
        n356) );
  MXI4X1 U2344 ( .A(\register[4][29] ), .B(\register[5][29] ), .C(
        \register[6][29] ), .D(\register[7][29] ), .S0(n494), .S1(n453), .Y(
        n376) );
  MXI4X1 U2345 ( .A(\register[20][29] ), .B(\register[21][29] ), .C(
        \register[22][29] ), .D(\register[23][29] ), .S0(n494), .S1(n453), .Y(
        n372) );
  MXI4X1 U2346 ( .A(\register[20][22] ), .B(\register[21][22] ), .C(
        \register[22][22] ), .D(\register[23][22] ), .S0(n489), .S1(n448), .Y(
        n315) );
  MXI4X1 U2347 ( .A(\register[4][22] ), .B(\register[5][22] ), .C(
        \register[6][22] ), .D(\register[7][22] ), .S0(n489), .S1(n448), .Y(
        n319) );
  MXI4X1 U2348 ( .A(\register[20][24] ), .B(\register[21][24] ), .C(
        \register[22][24] ), .D(\register[23][24] ), .S0(n490), .S1(n449), .Y(
        n331) );
  MXI4X1 U2349 ( .A(\register[4][24] ), .B(\register[5][24] ), .C(
        \register[6][24] ), .D(\register[7][24] ), .S0(n491), .S1(n450), .Y(
        n335) );
  MXI4X1 U2350 ( .A(\register[4][26] ), .B(\register[5][26] ), .C(
        \register[6][26] ), .D(\register[7][26] ), .S0(n492), .S1(n451), .Y(
        n352) );
  MXI4X1 U2351 ( .A(\register[20][26] ), .B(\register[21][26] ), .C(
        \register[22][26] ), .D(\register[23][26] ), .S0(n492), .S1(n451), .Y(
        n348) );
  MXI4X1 U2352 ( .A(\register[4][28] ), .B(\register[5][28] ), .C(
        \register[6][28] ), .D(\register[7][28] ), .S0(n493), .S1(n452), .Y(
        n368) );
  MXI4X1 U2353 ( .A(\register[20][28] ), .B(\register[21][28] ), .C(
        \register[22][28] ), .D(\register[23][28] ), .S0(n493), .S1(n452), .Y(
        n364) );
  MXI4X1 U2354 ( .A(\register[20][31] ), .B(\register[21][31] ), .C(
        \register[22][31] ), .D(\register[23][31] ), .S0(n495), .S1(n454), .Y(
        n388) );
  MXI4X1 U2355 ( .A(\register[4][31] ), .B(\register[5][31] ), .C(
        \register[6][31] ), .D(\register[7][31] ), .S0(n495), .S1(n454), .Y(
        n392) );
  MXI4X1 U2356 ( .A(\register[20][30] ), .B(\register[21][30] ), .C(
        \register[22][30] ), .D(\register[23][30] ), .S0(n494), .S1(n453), .Y(
        n380) );
  MXI4X1 U2357 ( .A(\register[4][30] ), .B(\register[5][30] ), .C(
        \register[6][30] ), .D(\register[7][30] ), .S0(n495), .S1(n454), .Y(
        n384) );
  MXI4X1 U2358 ( .A(\register[0][23] ), .B(\register[1][23] ), .C(
        \register[2][23] ), .D(\register[3][23] ), .S0(n490), .S1(n449), .Y(
        n328) );
  MXI4X1 U2359 ( .A(\register[16][25] ), .B(\register[17][25] ), .C(
        \register[18][25] ), .D(\register[19][25] ), .S0(n491), .S1(n450), .Y(
        n340) );
  MXI4X1 U2360 ( .A(\register[0][27] ), .B(\register[1][27] ), .C(
        \register[2][27] ), .D(\register[3][27] ), .S0(n493), .S1(n452), .Y(
        n361) );
  MXI4X1 U2361 ( .A(\register[16][27] ), .B(\register[17][27] ), .C(
        \register[18][27] ), .D(\register[19][27] ), .S0(n492), .S1(n451), .Y(
        n357) );
  MXI4X1 U2362 ( .A(\register[0][29] ), .B(\register[1][29] ), .C(
        \register[2][29] ), .D(\register[3][29] ), .S0(n494), .S1(n453), .Y(
        n377) );
  MXI4X1 U2363 ( .A(\register[16][29] ), .B(\register[17][29] ), .C(
        \register[18][29] ), .D(\register[19][29] ), .S0(n494), .S1(n453), .Y(
        n373) );
  MXI4X1 U2364 ( .A(\register[16][22] ), .B(\register[17][22] ), .C(
        \register[18][22] ), .D(\register[19][22] ), .S0(n489), .S1(n448), .Y(
        n316) );
  MXI4X1 U2365 ( .A(\register[16][24] ), .B(\register[17][24] ), .C(
        \register[18][24] ), .D(\register[19][24] ), .S0(n490), .S1(n449), .Y(
        n332) );
  MXI4X1 U2366 ( .A(\register[0][26] ), .B(\register[1][26] ), .C(
        \register[2][26] ), .D(\register[3][26] ), .S0(n492), .S1(n451), .Y(
        n353) );
  MXI4X1 U2367 ( .A(\register[16][26] ), .B(\register[17][26] ), .C(
        \register[18][26] ), .D(\register[19][26] ), .S0(n492), .S1(n451), .Y(
        n349) );
  MXI4X1 U2368 ( .A(\register[0][28] ), .B(\register[1][28] ), .C(
        \register[2][28] ), .D(\register[3][28] ), .S0(n493), .S1(n452), .Y(
        n369) );
  MXI4X1 U2369 ( .A(\register[16][28] ), .B(\register[17][28] ), .C(
        \register[18][28] ), .D(\register[19][28] ), .S0(n493), .S1(n452), .Y(
        n365) );
  MXI4X1 U2370 ( .A(\register[16][31] ), .B(\register[17][31] ), .C(
        \register[18][31] ), .D(\register[19][31] ), .S0(n495), .S1(n454), .Y(
        n389) );
  MXI4X1 U2371 ( .A(\register[16][30] ), .B(\register[17][30] ), .C(
        \register[18][30] ), .D(\register[19][30] ), .S0(n494), .S1(n453), .Y(
        n381) );
  MXI4X1 U2372 ( .A(\register[12][23] ), .B(\register[13][23] ), .C(
        \register[14][23] ), .D(\register[15][23] ), .S0(n490), .S1(n449), .Y(
        n325) );
  MXI4X1 U2373 ( .A(\register[28][23] ), .B(\register[29][23] ), .C(
        \register[30][23] ), .D(\register[31][23] ), .S0(n490), .S1(n449), .Y(
        n321) );
  MXI4X1 U2374 ( .A(\register[28][25] ), .B(\register[29][25] ), .C(
        \register[30][25] ), .D(\register[31][25] ), .S0(n491), .S1(n450), .Y(
        n337) );
  MXI4X1 U2375 ( .A(\register[12][25] ), .B(\register[13][25] ), .C(
        \register[14][25] ), .D(\register[15][25] ), .S0(n491), .S1(n450), .Y(
        n341) );
  MXI4X1 U2376 ( .A(\register[12][27] ), .B(\register[13][27] ), .C(
        \register[14][27] ), .D(\register[15][27] ), .S0(n493), .S1(n452), .Y(
        n358) );
  MXI4X1 U2377 ( .A(\register[12][29] ), .B(\register[13][29] ), .C(
        \register[14][29] ), .D(\register[15][29] ), .S0(n494), .S1(n453), .Y(
        n374) );
  MXI4X1 U2378 ( .A(\register[28][22] ), .B(\register[29][22] ), .C(
        \register[30][22] ), .D(\register[31][22] ), .S0(n489), .S1(n448), .Y(
        n313) );
  MXI4X1 U2379 ( .A(\register[12][22] ), .B(\register[13][22] ), .C(
        \register[14][22] ), .D(\register[15][22] ), .S0(n489), .S1(n448), .Y(
        n317) );
  MXI4X1 U2380 ( .A(\register[28][24] ), .B(\register[29][24] ), .C(
        \register[30][24] ), .D(\register[31][24] ), .S0(n490), .S1(n449), .Y(
        n329) );
  MXI4X1 U2381 ( .A(\register[12][24] ), .B(\register[13][24] ), .C(
        \register[14][24] ), .D(\register[15][24] ), .S0(n491), .S1(n450), .Y(
        n333) );
  MXI4X1 U2382 ( .A(\register[12][26] ), .B(\register[13][26] ), .C(
        \register[14][26] ), .D(\register[15][26] ), .S0(n492), .S1(n451), .Y(
        n350) );
  MXI4X1 U2383 ( .A(\register[12][28] ), .B(\register[13][28] ), .C(
        \register[14][28] ), .D(\register[15][28] ), .S0(n493), .S1(n452), .Y(
        n366) );
  MXI4X1 U2384 ( .A(\register[28][31] ), .B(\register[29][31] ), .C(
        \register[30][31] ), .D(\register[31][31] ), .S0(n495), .S1(n454), .Y(
        n386) );
  MXI4X1 U2385 ( .A(\register[12][31] ), .B(\register[13][31] ), .C(
        \register[14][31] ), .D(\register[15][31] ), .S0(n495), .S1(n454), .Y(
        n390) );
  MXI4X1 U2386 ( .A(\register[28][30] ), .B(\register[29][30] ), .C(
        \register[30][30] ), .D(\register[31][30] ), .S0(n494), .S1(n453), .Y(
        n378) );
  MXI4X1 U2387 ( .A(\register[12][30] ), .B(\register[13][30] ), .C(
        \register[14][30] ), .D(\register[15][30] ), .S0(n495), .S1(n454), .Y(
        n382) );
  MXI4X1 U2388 ( .A(\register[8][23] ), .B(\register[9][23] ), .C(
        \register[10][23] ), .D(\register[11][23] ), .S0(n490), .S1(n449), .Y(
        n326) );
  MXI4X1 U2389 ( .A(\register[24][23] ), .B(\register[25][23] ), .C(
        \register[26][23] ), .D(\register[27][23] ), .S0(n490), .S1(n449), .Y(
        n322) );
  MXI4X1 U2390 ( .A(\register[24][25] ), .B(\register[25][25] ), .C(
        \register[26][25] ), .D(\register[27][25] ), .S0(n491), .S1(n450), .Y(
        n338) );
  MXI4X1 U2391 ( .A(\register[8][25] ), .B(\register[9][25] ), .C(
        \register[10][25] ), .D(\register[11][25] ), .S0(n491), .S1(n450), .Y(
        n343) );
  MXI4X1 U2392 ( .A(\register[8][27] ), .B(\register[9][27] ), .C(
        \register[10][27] ), .D(\register[11][27] ), .S0(n493), .S1(n452), .Y(
        n359) );
  MXI4X1 U2393 ( .A(\register[24][27] ), .B(\register[25][27] ), .C(
        \register[26][27] ), .D(\register[27][27] ), .S0(n492), .S1(n451), .Y(
        n355) );
  MXI4X1 U2394 ( .A(\register[8][29] ), .B(\register[9][29] ), .C(
        \register[10][29] ), .D(\register[11][29] ), .S0(n494), .S1(n453), .Y(
        n375) );
  MXI4X1 U2395 ( .A(\register[24][29] ), .B(\register[25][29] ), .C(
        \register[26][29] ), .D(\register[27][29] ), .S0(n494), .S1(n453), .Y(
        n371) );
  MXI4X1 U2396 ( .A(\register[24][22] ), .B(\register[25][22] ), .C(
        \register[26][22] ), .D(\register[27][22] ), .S0(n489), .S1(n448), .Y(
        n314) );
  MXI4X1 U2397 ( .A(\register[8][22] ), .B(\register[9][22] ), .C(
        \register[10][22] ), .D(\register[11][22] ), .S0(n489), .S1(n448), .Y(
        n318) );
  MXI4X1 U2398 ( .A(\register[24][24] ), .B(\register[25][24] ), .C(
        \register[26][24] ), .D(\register[27][24] ), .S0(n490), .S1(n449), .Y(
        n330) );
  MXI4X1 U2399 ( .A(\register[8][24] ), .B(\register[9][24] ), .C(
        \register[10][24] ), .D(\register[11][24] ), .S0(n491), .S1(n450), .Y(
        n334) );
  MXI4X1 U2400 ( .A(\register[8][26] ), .B(\register[9][26] ), .C(
        \register[10][26] ), .D(\register[11][26] ), .S0(n492), .S1(n451), .Y(
        n351) );
  MXI4X1 U2401 ( .A(\register[24][26] ), .B(\register[25][26] ), .C(
        \register[26][26] ), .D(\register[27][26] ), .S0(n492), .S1(n451), .Y(
        n347) );
  MXI4X1 U2402 ( .A(\register[8][28] ), .B(\register[9][28] ), .C(
        \register[10][28] ), .D(\register[11][28] ), .S0(n493), .S1(n452), .Y(
        n367) );
  MXI4X1 U2403 ( .A(\register[24][28] ), .B(\register[25][28] ), .C(
        \register[26][28] ), .D(\register[27][28] ), .S0(n493), .S1(n452), .Y(
        n363) );
  MXI4X1 U2404 ( .A(\register[24][31] ), .B(\register[25][31] ), .C(
        \register[26][31] ), .D(\register[27][31] ), .S0(n495), .S1(n454), .Y(
        n387) );
  MXI4X1 U2405 ( .A(\register[8][31] ), .B(\register[9][31] ), .C(
        \register[10][31] ), .D(\register[11][31] ), .S0(n495), .S1(n454), .Y(
        n391) );
  MXI4X1 U2406 ( .A(\register[24][30] ), .B(\register[25][30] ), .C(
        \register[26][30] ), .D(\register[27][30] ), .S0(n494), .S1(n453), .Y(
        n379) );
  MXI4X1 U2407 ( .A(\register[8][30] ), .B(\register[9][30] ), .C(
        \register[10][30] ), .D(\register[11][30] ), .S0(n495), .S1(n454), .Y(
        n383) );
  CLKBUFX3 U2408 ( .A(n397), .Y(n394) );
  CLKBUFX3 U2409 ( .A(N471), .Y(n397) );
  CLKBUFX3 U2410 ( .A(n822), .Y(n819) );
  CLKBUFX3 U2411 ( .A(N476), .Y(n822) );
  CLKBUFX3 U2412 ( .A(n413), .Y(n408) );
  CLKBUFX3 U2413 ( .A(N469), .Y(n413) );
  CLKBUFX3 U2414 ( .A(N469), .Y(n414) );
  CLKBUFX3 U2415 ( .A(N469), .Y(n415) );
  CLKBUFX3 U2416 ( .A(N471), .Y(n398) );
  CLKBUFX3 U2417 ( .A(N476), .Y(n823) );
endmodule


module Sign_Extend ( data_i, data_o );
  input [15:0] data_i;
  output [31:0] data_o;
  wire   data_o_31, n1;
  assign data_o_31 = data_i[15];

  INVX1 U1 ( .A(n1), .Y(data_o[28]) );
  INVX1 U2 ( .A(n1), .Y(data_o[19]) );
  CLKINVX1 U3 ( .A(data_o[25]), .Y(n1) );
  CLKBUFX3 U4 ( .A(data_o_31), .Y(data_o[25]) );
  CLKBUFX3 U5 ( .A(data_o_31), .Y(data_o[30]) );
  CLKBUFX3 U6 ( .A(data_i[14]), .Y(data_o[14]) );
  CLKBUFX3 U7 ( .A(data_i[13]), .Y(data_o[13]) );
  CLKBUFX3 U8 ( .A(data_i[12]), .Y(data_o[12]) );
  CLKBUFX3 U9 ( .A(data_i[11]), .Y(data_o[11]) );
  CLKBUFX3 U10 ( .A(data_i[10]), .Y(data_o[10]) );
  CLKBUFX3 U11 ( .A(data_i[9]), .Y(data_o[9]) );
  CLKBUFX3 U12 ( .A(data_i[8]), .Y(data_o[8]) );
  CLKBUFX3 U13 ( .A(data_i[7]), .Y(data_o[7]) );
  CLKBUFX3 U14 ( .A(data_i[6]), .Y(data_o[6]) );
  CLKBUFX3 U15 ( .A(data_i[5]), .Y(data_o[5]) );
  CLKBUFX3 U16 ( .A(data_i[4]), .Y(data_o[4]) );
  CLKBUFX3 U17 ( .A(data_i[3]), .Y(data_o[3]) );
  CLKBUFX3 U18 ( .A(data_i[2]), .Y(data_o[2]) );
  CLKBUFX3 U19 ( .A(data_i[1]), .Y(data_o[1]) );
  CLKBUFX3 U20 ( .A(data_i[0]), .Y(data_o[0]) );
  CLKINVX1 U21 ( .A(n1), .Y(data_o[29]) );
  CLKINVX1 U22 ( .A(n1), .Y(data_o[27]) );
  CLKINVX1 U23 ( .A(n1), .Y(data_o[31]) );
  CLKINVX1 U24 ( .A(n1), .Y(data_o[24]) );
  CLKINVX1 U25 ( .A(n1), .Y(data_o[23]) );
  CLKINVX1 U26 ( .A(n1), .Y(data_o[22]) );
  CLKINVX1 U27 ( .A(n1), .Y(data_o[21]) );
  CLKINVX1 U28 ( .A(n1), .Y(data_o[20]) );
  CLKINVX1 U29 ( .A(n1), .Y(data_o[18]) );
  CLKINVX1 U30 ( .A(n1), .Y(data_o[17]) );
  CLKINVX1 U31 ( .A(n1), .Y(data_o[16]) );
  CLKINVX1 U32 ( .A(n1), .Y(data_o[15]) );
  CLKINVX1 U33 ( .A(n1), .Y(data_o[26]) );
endmodule


module MUX2_32b_0 ( data0_i, data1_i, sel_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  output [31:0] data_o;
  input sel_i;
  wire   n1, n2, n3, n4, n5;

  CLKMX2X2 U1 ( .A(data0_i[1]), .B(data1_i[1]), .S0(sel_i), .Y(data_o[1]) );
  CLKMX2X2 U2 ( .A(data0_i[2]), .B(data1_i[2]), .S0(sel_i), .Y(data_o[2]) );
  CLKMX2X3 U3 ( .A(data0_i[0]), .B(data1_i[0]), .S0(sel_i), .Y(data_o[0]) );
  CLKBUFX3 U4 ( .A(n5), .Y(n1) );
  CLKBUFX3 U5 ( .A(n5), .Y(n2) );
  CLKBUFX3 U6 ( .A(n5), .Y(n3) );
  CLKBUFX3 U7 ( .A(n5), .Y(n4) );
  AO22X1 U8 ( .A0(data1_i[8]), .A1(sel_i), .B0(data0_i[8]), .B1(n1), .Y(
        data_o[8]) );
  AO22X1 U9 ( .A0(data1_i[3]), .A1(sel_i), .B0(data0_i[3]), .B1(n3), .Y(
        data_o[3]) );
  AO22X1 U10 ( .A0(data1_i[4]), .A1(sel_i), .B0(data0_i[4]), .B1(n3), .Y(
        data_o[4]) );
  AO22X1 U11 ( .A0(data1_i[5]), .A1(sel_i), .B0(data0_i[5]), .B1(n3), .Y(
        data_o[5]) );
  AO22X1 U12 ( .A0(data1_i[6]), .A1(sel_i), .B0(data0_i[6]), .B1(n2), .Y(
        data_o[6]) );
  AO22X1 U13 ( .A0(data1_i[7]), .A1(sel_i), .B0(data0_i[7]), .B1(n2), .Y(
        data_o[7]) );
  AO22X1 U14 ( .A0(data1_i[10]), .A1(sel_i), .B0(data0_i[10]), .B1(n4), .Y(
        data_o[10]) );
  AO22X1 U15 ( .A0(sel_i), .A1(data1_i[9]), .B0(data0_i[9]), .B1(n1), .Y(
        data_o[9]) );
  AO22X1 U16 ( .A0(data1_i[18]), .A1(sel_i), .B0(data0_i[18]), .B1(n3), .Y(
        data_o[18]) );
  AO22X1 U17 ( .A0(data1_i[11]), .A1(sel_i), .B0(data0_i[11]), .B1(n4), .Y(
        data_o[11]) );
  AO22X1 U18 ( .A0(data1_i[12]), .A1(sel_i), .B0(data0_i[12]), .B1(n4), .Y(
        data_o[12]) );
  AO22X1 U19 ( .A0(data1_i[13]), .A1(sel_i), .B0(data0_i[13]), .B1(n4), .Y(
        data_o[13]) );
  AO22X1 U20 ( .A0(data1_i[19]), .A1(sel_i), .B0(data0_i[19]), .B1(n3), .Y(
        data_o[19]) );
  AO22X1 U21 ( .A0(data1_i[20]), .A1(sel_i), .B0(data0_i[20]), .B1(n3), .Y(
        data_o[20]) );
  AO22X1 U22 ( .A0(data1_i[21]), .A1(sel_i), .B0(data0_i[21]), .B1(n3), .Y(
        data_o[21]) );
  AO22X1 U23 ( .A0(data1_i[15]), .A1(sel_i), .B0(data0_i[15]), .B1(n4), .Y(
        data_o[15]) );
  AO22X1 U24 ( .A0(data1_i[16]), .A1(sel_i), .B0(data0_i[16]), .B1(n4), .Y(
        data_o[16]) );
  AO22X1 U25 ( .A0(data1_i[17]), .A1(sel_i), .B0(data0_i[17]), .B1(n4), .Y(
        data_o[17]) );
  AO22X1 U26 ( .A0(data1_i[14]), .A1(sel_i), .B0(data0_i[14]), .B1(n4), .Y(
        data_o[14]) );
  AO22X1 U27 ( .A0(data1_i[22]), .A1(sel_i), .B0(data0_i[22]), .B1(n3), .Y(
        data_o[22]) );
  AO22X1 U28 ( .A0(data1_i[26]), .A1(sel_i), .B0(data0_i[26]), .B1(n3), .Y(
        data_o[26]) );
  AO22X1 U29 ( .A0(data1_i[27]), .A1(sel_i), .B0(data0_i[27]), .B1(n3), .Y(
        data_o[27]) );
  AO22X1 U30 ( .A0(data1_i[28]), .A1(sel_i), .B0(data0_i[28]), .B1(n3), .Y(
        data_o[28]) );
  AO22X1 U31 ( .A0(data1_i[29]), .A1(sel_i), .B0(data0_i[29]), .B1(n3), .Y(
        data_o[29]) );
  AO22X1 U32 ( .A0(data1_i[23]), .A1(sel_i), .B0(data0_i[23]), .B1(n3), .Y(
        data_o[23]) );
  AO22X1 U33 ( .A0(data1_i[24]), .A1(sel_i), .B0(data0_i[24]), .B1(n3), .Y(
        data_o[24]) );
  AO22X1 U34 ( .A0(data1_i[25]), .A1(sel_i), .B0(data0_i[25]), .B1(n3), .Y(
        data_o[25]) );
  AO22X1 U35 ( .A0(data1_i[30]), .A1(sel_i), .B0(data0_i[30]), .B1(n3), .Y(
        data_o[30]) );
  AO22X1 U36 ( .A0(data1_i[31]), .A1(sel_i), .B0(data0_i[31]), .B1(n3), .Y(
        data_o[31]) );
  CLKINVX1 U37 ( .A(sel_i), .Y(n5) );
endmodule


module ALU_Control ( func_i, ALUOp_i, ALUctrl_o );
  input [3:0] func_i;
  input [1:0] ALUOp_i;
  output [2:0] ALUctrl_o;
  wire   n5, n6, n7, n8, n1, n2, n3, n4;

  CLKINVX1 U3 ( .A(ALUOp_i[0]), .Y(n1) );
  NAND3X1 U4 ( .A(ALUOp_i[1]), .B(n1), .C(n7), .Y(n5) );
  NOR2X1 U5 ( .A(n8), .B(n5), .Y(ALUctrl_o[0]) );
  AOI33X1 U6 ( .A0(func_i[1]), .A1(n4), .A2(func_i[3]), .B0(n3), .B1(n2), .B2(
        func_i[0]), .Y(n8) );
  OAI32X1 U7 ( .A0(n3), .A1(func_i[0]), .A2(n5), .B0(ALUOp_i[1]), .B1(n1), .Y(
        ALUctrl_o[2]) );
  OAI31XL U8 ( .A0(n6), .A1(func_i[0]), .A2(ALUOp_i[0]), .B0(ALUOp_i[1]), .Y(
        ALUctrl_o[1]) );
  OAI21XL U9 ( .A0(func_i[1]), .A1(n2), .B0(n7), .Y(n6) );
  XOR2X1 U10 ( .A(n4), .B(func_i[2]), .Y(n7) );
  CLKINVX1 U11 ( .A(func_i[0]), .Y(n4) );
  CLKINVX1 U12 ( .A(func_i[3]), .Y(n2) );
  CLKINVX1 U13 ( .A(func_i[1]), .Y(n3) );
endmodule


module ALU_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104;

  INVXL U1 ( .A(A[1]), .Y(n30) );
  NOR2XL U2 ( .A(n25), .B(B[6]), .Y(n99) );
  NOR2XL U3 ( .A(n27), .B(B[4]), .Y(n104) );
  INVXL U4 ( .A(B[3]), .Y(n28) );
  NOR2BXL U5 ( .AN(A[5]), .B(B[5]), .Y(n98) );
  NAND2XL U6 ( .A(A[3]), .B(n28), .Y(n60) );
  NAND2XL U7 ( .A(A[2]), .B(n29), .Y(n59) );
  NAND2BXL U8 ( .AN(A[5]), .B(B[5]), .Y(n97) );
  INVXL U9 ( .A(B[1]), .Y(n31) );
  NOR2BXL U10 ( .AN(A[0]), .B(B[0]), .Y(n40) );
  CLKINVX1 U11 ( .A(B[2]), .Y(n29) );
  CLKINVX1 U12 ( .A(B[9]), .Y(n22) );
  CLKINVX1 U13 ( .A(B[10]), .Y(n21) );
  CLKINVX1 U14 ( .A(B[19]), .Y(n13) );
  CLKINVX1 U15 ( .A(B[11]), .Y(n20) );
  CLKINVX1 U16 ( .A(B[13]), .Y(n18) );
  CLKINVX1 U17 ( .A(B[21]), .Y(n11) );
  CLKINVX1 U18 ( .A(B[12]), .Y(n19) );
  CLKINVX1 U19 ( .A(B[20]), .Y(n12) );
  CLKINVX1 U20 ( .A(B[18]), .Y(n14) );
  CLKINVX1 U21 ( .A(B[26]), .Y(n7) );
  CLKINVX1 U22 ( .A(B[27]), .Y(n5) );
  CLKINVX1 U23 ( .A(B[29]), .Y(n3) );
  CLKINVX1 U24 ( .A(B[28]), .Y(n4) );
  CLKINVX1 U25 ( .A(A[31]), .Y(n1) );
  CLKINVX1 U26 ( .A(B[8]), .Y(n23) );
  CLKINVX1 U27 ( .A(n104), .Y(n26) );
  CLKINVX1 U28 ( .A(n44), .Y(n6) );
  CLKINVX1 U29 ( .A(A[4]), .Y(n27) );
  CLKINVX1 U30 ( .A(A[7]), .Y(n24) );
  CLKINVX1 U31 ( .A(A[6]), .Y(n25) );
  CLKINVX1 U32 ( .A(A[17]), .Y(n15) );
  CLKINVX1 U33 ( .A(A[16]), .Y(n16) );
  CLKINVX1 U34 ( .A(A[14]), .Y(n17) );
  CLKINVX1 U35 ( .A(A[25]), .Y(n8) );
  CLKINVX1 U36 ( .A(A[24]), .Y(n9) );
  CLKINVX1 U37 ( .A(A[22]), .Y(n10) );
  CLKINVX1 U38 ( .A(A[30]), .Y(n2) );
  NOR4X1 U39 ( .A(n32), .B(n33), .C(n34), .D(n35), .Y(EQ) );
  NAND4X1 U40 ( .A(n36), .B(n37), .C(n38), .D(n39), .Y(n35) );
  OAI22XL U41 ( .A0(A[1]), .A1(n40), .B0(n40), .B1(n31), .Y(n36) );
  NAND4BBXL U42 ( .AN(n41), .BN(n42), .C(n43), .D(n44), .Y(n34) );
  NAND2BX1 U43 ( .AN(n45), .B(n46), .Y(n33) );
  NOR4BX1 U44 ( .AN(n47), .B(n48), .C(n49), .D(n50), .Y(n46) );
  NAND4BX1 U45 ( .AN(n51), .B(n52), .C(n53), .D(n54), .Y(n45) );
  NAND4BBXL U46 ( .AN(n55), .BN(n56), .C(n57), .D(n58), .Y(n32) );
  NOR4BBX1 U47 ( .AN(n59), .BN(n60), .C(LT), .D(n61), .Y(n58) );
  OAI22XL U48 ( .A0(B[31]), .A1(n1), .B0(n61), .B1(n62), .Y(LT) );
  AOI32X1 U49 ( .A0(n37), .A1(n38), .A2(n63), .B0(B[30]), .B1(n2), .Y(n62) );
  OAI221XL U50 ( .A0(A[28]), .A1(n4), .B0(A[29]), .B1(n3), .C0(n64), .Y(n63)
         );
  OAI211X1 U51 ( .A0(n65), .A1(n66), .B0(n39), .C0(n43), .Y(n64) );
  NAND2X1 U52 ( .A(A[27]), .B(n5), .Y(n43) );
  NAND2X1 U53 ( .A(A[28]), .B(n4), .Y(n39) );
  OAI32X1 U54 ( .A0(n67), .A1(n41), .A2(n6), .B0(A[26]), .B1(n7), .Y(n66) );
  NAND2X1 U55 ( .A(A[26]), .B(n7), .Y(n44) );
  NOR2X1 U56 ( .A(n8), .B(B[25]), .Y(n41) );
  AOI221XL U57 ( .A0(B[25]), .A1(n8), .B0(B[24]), .B1(n9), .C0(n68), .Y(n67)
         );
  AOI211X1 U58 ( .A0(n69), .A1(n70), .B0(n51), .C0(n42), .Y(n68) );
  NOR2X1 U59 ( .A(n9), .B(B[24]), .Y(n42) );
  NOR2BX1 U60 ( .AN(A[23]), .B(B[23]), .Y(n51) );
  NAND2BX1 U61 ( .AN(A[23]), .B(B[23]), .Y(n70) );
  AOI32X1 U62 ( .A0(n54), .A1(n53), .A2(n71), .B0(B[22]), .B1(n10), .Y(n69) );
  OAI221XL U63 ( .A0(A[20]), .A1(n12), .B0(A[21]), .B1(n11), .C0(n72), .Y(n71)
         );
  OAI211X1 U64 ( .A0(n73), .A1(n74), .B0(n52), .C0(n47), .Y(n72) );
  NAND2X1 U65 ( .A(A[19]), .B(n13), .Y(n47) );
  NAND2X1 U66 ( .A(A[20]), .B(n12), .Y(n52) );
  OAI32X1 U67 ( .A0(n75), .A1(n49), .A2(n50), .B0(A[18]), .B1(n14), .Y(n74) );
  NOR2BX1 U68 ( .AN(A[18]), .B(B[18]), .Y(n50) );
  NOR2X1 U69 ( .A(n15), .B(B[17]), .Y(n49) );
  AOI221XL U70 ( .A0(B[17]), .A1(n15), .B0(B[16]), .B1(n16), .C0(n76), .Y(n75)
         );
  AOI211X1 U71 ( .A0(n77), .A1(n78), .B0(n79), .C0(n48), .Y(n76) );
  NOR2X1 U72 ( .A(n16), .B(B[16]), .Y(n48) );
  NAND2BX1 U73 ( .AN(A[15]), .B(B[15]), .Y(n78) );
  AOI32X1 U74 ( .A0(n80), .A1(n81), .A2(n82), .B0(B[14]), .B1(n17), .Y(n77) );
  OAI221XL U75 ( .A0(A[12]), .A1(n19), .B0(A[13]), .B1(n18), .C0(n83), .Y(n82)
         );
  NAND3X1 U76 ( .A(n84), .B(n85), .C(n86), .Y(n83) );
  OAI221XL U77 ( .A0(A[10]), .A1(n21), .B0(A[11]), .B1(n20), .C0(n87), .Y(n86)
         );
  OAI211X1 U78 ( .A0(n88), .A1(n89), .B0(n90), .C0(n91), .Y(n87) );
  OAI32X1 U79 ( .A0(n92), .A1(n93), .A2(n94), .B0(A[8]), .B1(n23), .Y(n89) );
  AOI221XL U80 ( .A0(B[7]), .A1(n24), .B0(B[6]), .B1(n25), .C0(n95), .Y(n92)
         );
  AOI211X1 U81 ( .A0(n96), .A1(n97), .B0(n98), .C0(n99), .Y(n95) );
  AOI32X1 U82 ( .A0(n26), .A1(n60), .A2(n100), .B0(B[4]), .B1(n27), .Y(n96) );
  OAI221XL U83 ( .A0(A[2]), .A1(n29), .B0(A[3]), .B1(n28), .C0(n101), .Y(n100)
         );
  OAI211X1 U84 ( .A0(n102), .A1(n30), .B0(n103), .C0(n59), .Y(n101) );
  AO21X1 U85 ( .A0(n30), .A1(n102), .B0(B[1]), .Y(n103) );
  NOR2BX1 U86 ( .AN(B[0]), .B(A[0]), .Y(n102) );
  NOR2X1 U87 ( .A(A[9]), .B(n22), .Y(n88) );
  NOR2X1 U88 ( .A(A[19]), .B(n13), .Y(n73) );
  NAND2X1 U89 ( .A(A[21]), .B(n11), .Y(n53) );
  NAND2BX1 U90 ( .AN(B[22]), .B(A[22]), .Y(n54) );
  NOR2X1 U91 ( .A(A[27]), .B(n5), .Y(n65) );
  OR2X1 U92 ( .A(B[30]), .B(n2), .Y(n38) );
  NAND2X1 U93 ( .A(A[29]), .B(n3), .Y(n37) );
  NOR2BX1 U94 ( .AN(B[31]), .B(A[31]), .Y(n61) );
  NOR4X1 U95 ( .A(n104), .B(n98), .C(n99), .D(n93), .Y(n57) );
  NOR2X1 U96 ( .A(n24), .B(B[7]), .Y(n93) );
  NAND4BX1 U97 ( .AN(n94), .B(n91), .C(n90), .D(n85), .Y(n56) );
  NAND2X1 U98 ( .A(A[11]), .B(n20), .Y(n85) );
  NAND2X1 U99 ( .A(A[10]), .B(n21), .Y(n90) );
  NAND2X1 U100 ( .A(A[9]), .B(n22), .Y(n91) );
  NOR2BX1 U101 ( .AN(A[8]), .B(B[8]), .Y(n94) );
  NAND4BX1 U102 ( .AN(n79), .B(n84), .C(n81), .D(n80), .Y(n55) );
  NAND2BX1 U103 ( .AN(B[14]), .B(A[14]), .Y(n80) );
  NAND2X1 U104 ( .A(A[13]), .B(n18), .Y(n81) );
  NAND2X1 U105 ( .A(A[12]), .B(n19), .Y(n84) );
  NOR2BX1 U106 ( .AN(A[15]), .B(B[15]), .Y(n79) );
endmodule


module ALU_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n37, n39, n40, n41, n42, n43, n45, n47, n48,
         n49, n50, n51, n53, n55, n56, n57, n58, n59, n61, n63, n64, n65, n66,
         n67, n69, n71, n72, n73, n74, n75, n77, n79, n80, n81, n82, n83, n85,
         n87, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99, n101, n103,
         n104, n105, n106, n107, n109, n111, n112, n113, n114, n115, n117,
         n119, n120, n121, n122, n123, n125, n127, n128, n129, n130, n132,
         n134, n135, n137, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n180, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330;

  ADDFXL U3 ( .A(n184), .B(A[30]), .CI(n32), .CO(n31), .S(DIFF[30]) );
  XOR2X1 U4 ( .A(n35), .B(n2), .Y(DIFF[29]) );
  XOR2X1 U18 ( .A(n43), .B(n4), .Y(DIFF[27]) );
  XOR2X1 U32 ( .A(n51), .B(n6), .Y(DIFF[25]) );
  XOR2X1 U46 ( .A(n59), .B(n8), .Y(DIFF[23]) );
  XOR2X1 U60 ( .A(n67), .B(n10), .Y(DIFF[21]) );
  XOR2X1 U74 ( .A(n75), .B(n12), .Y(DIFF[19]) );
  XOR2X1 U88 ( .A(n83), .B(n14), .Y(DIFF[17]) );
  XOR2X1 U102 ( .A(n91), .B(n16), .Y(DIFF[15]) );
  XOR2X1 U116 ( .A(n99), .B(n18), .Y(DIFF[13]) );
  XOR2X1 U130 ( .A(n107), .B(n20), .Y(DIFF[11]) );
  XOR2X1 U144 ( .A(n115), .B(n22), .Y(DIFF[9]) );
  XOR2X1 U158 ( .A(n123), .B(n24), .Y(DIFF[7]) );
  XOR2X1 U172 ( .A(n135), .B(n26), .Y(DIFF[5]) );
  XOR2X1 U199 ( .A(n149), .B(n29), .Y(DIFF[2]) );
  XOR2X1 U205 ( .A(n30), .B(n153), .Y(DIFF[1]) );
  XNOR2XL U249 ( .A(n128), .B(n25), .Y(DIFF[6]) );
  NOR2XL U250 ( .A(n213), .B(A[1]), .Y(n151) );
  OAI21XL U251 ( .A0(n141), .A1(n129), .B0(n130), .Y(n128) );
  OAI21X1 U252 ( .A0(n123), .A1(n121), .B0(n122), .Y(n120) );
  OAI21XL U253 ( .A0(n35), .A1(n33), .B0(n34), .Y(n32) );
  NAND2BX1 U254 ( .AN(n147), .B(n148), .Y(n29) );
  NAND2BX1 U255 ( .AN(n121), .B(n122), .Y(n24) );
  AOI21XL U256 ( .A0(n140), .A1(n317), .B0(n137), .Y(n135) );
  NAND2XL U257 ( .A(n318), .B(n134), .Y(n26) );
  XNOR2XL U258 ( .A(n120), .B(n23), .Y(DIFF[8]) );
  NAND2XL U259 ( .A(n317), .B(n139), .Y(n27) );
  AOI21XL U260 ( .A0(n128), .A1(n319), .B0(n125), .Y(n123) );
  AOI21XL U261 ( .A0(n120), .A1(n320), .B0(n117), .Y(n115) );
  AOI21XL U262 ( .A0(n112), .A1(n323), .B0(n109), .Y(n107) );
  AOI21XL U263 ( .A0(n104), .A1(n324), .B0(n101), .Y(n99) );
  AOI21XL U264 ( .A0(n96), .A1(n321), .B0(n93), .Y(n91) );
  AOI21XL U265 ( .A0(n88), .A1(n322), .B0(n85), .Y(n83) );
  AOI21XL U266 ( .A0(n80), .A1(n326), .B0(n77), .Y(n75) );
  AOI21XL U267 ( .A0(n72), .A1(n325), .B0(n69), .Y(n67) );
  AOI21XL U268 ( .A0(n64), .A1(n328), .B0(n61), .Y(n59) );
  AOI21XL U269 ( .A0(n56), .A1(n327), .B0(n53), .Y(n51) );
  AOI21XL U270 ( .A0(n48), .A1(n329), .B0(n45), .Y(n43) );
  AOI21XL U271 ( .A0(n40), .A1(n330), .B0(n37), .Y(n35) );
  AOI21XL U272 ( .A0(n150), .A1(n142), .B0(n143), .Y(n141) );
  OAI21X1 U273 ( .A0(n148), .A1(n144), .B0(n145), .Y(n143) );
  XNOR2XL U274 ( .A(n40), .B(n3), .Y(DIFF[28]) );
  XNOR2XL U275 ( .A(n64), .B(n9), .Y(DIFF[22]) );
  XNOR2XL U276 ( .A(n56), .B(n7), .Y(DIFF[24]) );
  XNOR2XL U277 ( .A(n48), .B(n5), .Y(DIFF[26]) );
  XNOR2XL U278 ( .A(n80), .B(n13), .Y(DIFF[18]) );
  XNOR2XL U279 ( .A(n96), .B(n17), .Y(DIFF[14]) );
  XNOR2XL U280 ( .A(n88), .B(n15), .Y(DIFF[16]) );
  XNOR2XL U281 ( .A(n72), .B(n11), .Y(DIFF[20]) );
  XNOR2XL U282 ( .A(n112), .B(n21), .Y(DIFF[10]) );
  XNOR2XL U283 ( .A(n104), .B(n19), .Y(DIFF[12]) );
  NAND2BXL U284 ( .AN(n151), .B(n152), .Y(n30) );
  NAND2XL U285 ( .A(n208), .B(A[6]), .Y(n127) );
  NAND2XL U286 ( .A(n209), .B(A[5]), .Y(n134) );
  NAND2XL U287 ( .A(n210), .B(A[4]), .Y(n139) );
  NOR2XL U288 ( .A(n212), .B(A[2]), .Y(n147) );
  NOR2X1 U289 ( .A(n211), .B(A[3]), .Y(n144) );
  NAND2XL U290 ( .A(n211), .B(A[3]), .Y(n145) );
  NAND2XL U291 ( .A(n213), .B(A[1]), .Y(n152) );
  XOR2XL U292 ( .A(n31), .B(n1), .Y(DIFF[31]) );
  XNOR2XL U293 ( .A(n214), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U294 ( .A(n141), .Y(n140) );
  CLKINVX1 U295 ( .A(n150), .Y(n149) );
  OAI21XL U296 ( .A0(n151), .A1(n153), .B0(n152), .Y(n150) );
  NOR2X1 U297 ( .A(n147), .B(n144), .Y(n142) );
  AOI21X1 U298 ( .A0(n318), .A1(n137), .B0(n132), .Y(n130) );
  NAND2X1 U299 ( .A(n317), .B(n318), .Y(n129) );
  CLKINVX1 U300 ( .A(n134), .Y(n132) );
  NAND2X1 U301 ( .A(n320), .B(n119), .Y(n23) );
  XNOR2X1 U302 ( .A(n146), .B(n28), .Y(DIFF[3]) );
  NAND2X1 U303 ( .A(n180), .B(n145), .Y(n28) );
  OAI21XL U304 ( .A0(n149), .A1(n147), .B0(n148), .Y(n146) );
  CLKINVX1 U305 ( .A(n144), .Y(n180) );
  XNOR2X1 U306 ( .A(n140), .B(n27), .Y(DIFF[4]) );
  NAND2X1 U307 ( .A(n319), .B(n127), .Y(n25) );
  CLKINVX1 U308 ( .A(n127), .Y(n125) );
  CLKINVX1 U309 ( .A(B[1]), .Y(n213) );
  CLKINVX1 U310 ( .A(B[2]), .Y(n212) );
  CLKINVX1 U311 ( .A(B[8]), .Y(n206) );
  CLKINVX1 U312 ( .A(B[3]), .Y(n211) );
  CLKINVX1 U313 ( .A(B[4]), .Y(n210) );
  CLKINVX1 U314 ( .A(B[5]), .Y(n209) );
  CLKINVX1 U315 ( .A(B[6]), .Y(n208) );
  CLKINVX1 U316 ( .A(B[7]), .Y(n207) );
  CLKINVX1 U317 ( .A(B[0]), .Y(n214) );
  CLKINVX1 U318 ( .A(n139), .Y(n137) );
  OAI21XL U319 ( .A0(n83), .A1(n81), .B0(n82), .Y(n80) );
  OAI21XL U320 ( .A0(n51), .A1(n49), .B0(n50), .Y(n48) );
  OAI21XL U321 ( .A0(n115), .A1(n113), .B0(n114), .Y(n112) );
  OAI21XL U322 ( .A0(n75), .A1(n73), .B0(n74), .Y(n72) );
  OAI21XL U323 ( .A0(n43), .A1(n41), .B0(n42), .Y(n40) );
  OAI21XL U324 ( .A0(n107), .A1(n105), .B0(n106), .Y(n104) );
  OAI21XL U325 ( .A0(n99), .A1(n97), .B0(n98), .Y(n96) );
  OAI21XL U326 ( .A0(n67), .A1(n65), .B0(n66), .Y(n64) );
  OAI21XL U327 ( .A0(n91), .A1(n89), .B0(n90), .Y(n88) );
  OAI21XL U328 ( .A0(n59), .A1(n57), .B0(n58), .Y(n56) );
  CLKINVX1 U329 ( .A(n119), .Y(n117) );
  CLKINVX1 U330 ( .A(n111), .Y(n109) );
  CLKINVX1 U331 ( .A(n103), .Y(n101) );
  CLKINVX1 U332 ( .A(n95), .Y(n93) );
  CLKINVX1 U333 ( .A(n87), .Y(n85) );
  CLKINVX1 U334 ( .A(n79), .Y(n77) );
  CLKINVX1 U335 ( .A(n71), .Y(n69) );
  CLKINVX1 U336 ( .A(n63), .Y(n61) );
  CLKINVX1 U337 ( .A(n55), .Y(n53) );
  CLKINVX1 U338 ( .A(n47), .Y(n45) );
  CLKINVX1 U339 ( .A(n39), .Y(n37) );
  CLKINVX1 U340 ( .A(B[18]), .Y(n196) );
  CLKINVX1 U341 ( .A(B[11]), .Y(n203) );
  CLKINVX1 U342 ( .A(B[13]), .Y(n201) );
  CLKINVX1 U343 ( .A(B[19]), .Y(n195) );
  CLKINVX1 U344 ( .A(B[21]), .Y(n193) );
  CLKINVX1 U345 ( .A(B[10]), .Y(n204) );
  CLKINVX1 U346 ( .A(B[12]), .Y(n202) );
  CLKINVX1 U347 ( .A(B[20]), .Y(n194) );
  CLKINVX1 U348 ( .A(B[9]), .Y(n205) );
  CLKINVX1 U349 ( .A(B[15]), .Y(n199) );
  CLKINVX1 U350 ( .A(B[16]), .Y(n198) );
  CLKINVX1 U351 ( .A(B[17]), .Y(n197) );
  CLKINVX1 U352 ( .A(B[14]), .Y(n200) );
  CLKINVX1 U353 ( .A(B[27]), .Y(n187) );
  CLKINVX1 U354 ( .A(B[29]), .Y(n185) );
  CLKINVX1 U355 ( .A(B[26]), .Y(n188) );
  CLKINVX1 U356 ( .A(B[28]), .Y(n186) );
  CLKINVX1 U357 ( .A(B[23]), .Y(n191) );
  CLKINVX1 U358 ( .A(B[24]), .Y(n190) );
  CLKINVX1 U359 ( .A(B[25]), .Y(n189) );
  CLKINVX1 U360 ( .A(B[22]), .Y(n192) );
  NAND2X1 U361 ( .A(n321), .B(n95), .Y(n17) );
  NAND2X1 U362 ( .A(n328), .B(n63), .Y(n9) );
  NAND2X1 U363 ( .A(n322), .B(n87), .Y(n15) );
  NAND2X1 U364 ( .A(n327), .B(n55), .Y(n7) );
  NAND2X1 U365 ( .A(n329), .B(n47), .Y(n5) );
  NAND2X1 U366 ( .A(n323), .B(n111), .Y(n21) );
  NAND2X1 U367 ( .A(n324), .B(n103), .Y(n19) );
  NAND2X1 U368 ( .A(n325), .B(n71), .Y(n11) );
  NAND2X1 U369 ( .A(n330), .B(n39), .Y(n3) );
  NAND2X1 U370 ( .A(n326), .B(n79), .Y(n13) );
  NAND2BX1 U371 ( .AN(n113), .B(n114), .Y(n22) );
  NAND2BX1 U372 ( .AN(n81), .B(n82), .Y(n14) );
  NAND2BX1 U373 ( .AN(n49), .B(n50), .Y(n6) );
  NAND2BX1 U374 ( .AN(n73), .B(n74), .Y(n12) );
  NAND2BX1 U375 ( .AN(n41), .B(n42), .Y(n4) );
  NAND2BX1 U376 ( .AN(n105), .B(n106), .Y(n20) );
  NAND2BX1 U377 ( .AN(n97), .B(n98), .Y(n18) );
  NAND2BX1 U378 ( .AN(n65), .B(n66), .Y(n10) );
  NAND2BX1 U379 ( .AN(n33), .B(n34), .Y(n2) );
  NAND2BX1 U380 ( .AN(n89), .B(n90), .Y(n16) );
  NAND2BX1 U381 ( .AN(n57), .B(n58), .Y(n8) );
  NAND2X1 U382 ( .A(n212), .B(A[2]), .Y(n148) );
  NOR2X1 U383 ( .A(n207), .B(A[7]), .Y(n121) );
  NAND2X1 U384 ( .A(n207), .B(A[7]), .Y(n122) );
  NAND2X1 U385 ( .A(n206), .B(A[8]), .Y(n119) );
  NOR2X1 U386 ( .A(n214), .B(A[0]), .Y(n153) );
  OR2X1 U387 ( .A(n210), .B(A[4]), .Y(n317) );
  OR2X1 U388 ( .A(n209), .B(A[5]), .Y(n318) );
  OR2X1 U389 ( .A(n208), .B(A[6]), .Y(n319) );
  OR2X1 U390 ( .A(n206), .B(A[8]), .Y(n320) );
  CLKINVX1 U391 ( .A(B[30]), .Y(n184) );
  NAND2X1 U392 ( .A(n200), .B(A[14]), .Y(n95) );
  NOR2X1 U393 ( .A(n197), .B(A[17]), .Y(n81) );
  NAND2X1 U394 ( .A(n198), .B(A[16]), .Y(n87) );
  NOR2X1 U395 ( .A(n205), .B(A[9]), .Y(n113) );
  NOR2X1 U396 ( .A(n195), .B(A[19]), .Y(n73) );
  NAND2X1 U397 ( .A(n197), .B(A[17]), .Y(n82) );
  NOR2X1 U398 ( .A(n203), .B(A[11]), .Y(n105) );
  NOR2X1 U399 ( .A(n201), .B(A[13]), .Y(n97) );
  NOR2X1 U400 ( .A(n193), .B(A[21]), .Y(n65) );
  NAND2X1 U401 ( .A(n204), .B(A[10]), .Y(n111) );
  NAND2X1 U402 ( .A(n202), .B(A[12]), .Y(n103) );
  NAND2X1 U403 ( .A(n194), .B(A[20]), .Y(n71) );
  NAND2X1 U404 ( .A(n196), .B(A[18]), .Y(n79) );
  NOR2X1 U405 ( .A(n199), .B(A[15]), .Y(n89) );
  NAND2X1 U406 ( .A(n205), .B(A[9]), .Y(n114) );
  NAND2X1 U407 ( .A(n195), .B(A[19]), .Y(n74) );
  NAND2X1 U408 ( .A(n203), .B(A[11]), .Y(n106) );
  NAND2X1 U409 ( .A(n201), .B(A[13]), .Y(n98) );
  NAND2X1 U410 ( .A(n199), .B(A[15]), .Y(n90) );
  OR2X1 U411 ( .A(n200), .B(A[14]), .Y(n321) );
  OR2X1 U412 ( .A(n198), .B(A[16]), .Y(n322) );
  OR2X1 U413 ( .A(n204), .B(A[10]), .Y(n323) );
  OR2X1 U414 ( .A(n202), .B(A[12]), .Y(n324) );
  OR2X1 U415 ( .A(n194), .B(A[20]), .Y(n325) );
  OR2X1 U416 ( .A(n196), .B(A[18]), .Y(n326) );
  XNOR2X1 U417 ( .A(B[31]), .B(A[31]), .Y(n1) );
  NAND2X1 U418 ( .A(n192), .B(A[22]), .Y(n63) );
  NOR2X1 U419 ( .A(n189), .B(A[25]), .Y(n49) );
  NAND2X1 U420 ( .A(n190), .B(A[24]), .Y(n55) );
  NOR2X1 U421 ( .A(n187), .B(A[27]), .Y(n41) );
  NAND2X1 U422 ( .A(n189), .B(A[25]), .Y(n50) );
  NOR2X1 U423 ( .A(n185), .B(A[29]), .Y(n33) );
  NAND2X1 U424 ( .A(n188), .B(A[26]), .Y(n47) );
  NAND2X1 U425 ( .A(n186), .B(A[28]), .Y(n39) );
  NOR2X1 U426 ( .A(n191), .B(A[23]), .Y(n57) );
  NAND2X1 U427 ( .A(n187), .B(A[27]), .Y(n42) );
  NAND2X1 U428 ( .A(n193), .B(A[21]), .Y(n66) );
  NAND2X1 U429 ( .A(n185), .B(A[29]), .Y(n34) );
  NAND2X1 U430 ( .A(n191), .B(A[23]), .Y(n58) );
  OR2X1 U431 ( .A(n190), .B(A[24]), .Y(n327) );
  OR2X1 U432 ( .A(n192), .B(A[22]), .Y(n328) );
  OR2X1 U433 ( .A(n188), .B(A[26]), .Y(n329) );
  OR2X1 U434 ( .A(n186), .B(A[28]), .Y(n330) );
endmodule


module ALU_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n38, n40, n41, n42, n43, n44, n46, n48,
         n49, n50, n51, n52, n54, n56, n57, n58, n59, n60, n62, n64, n65, n66,
         n67, n68, n70, n72, n73, n74, n75, n76, n78, n80, n81, n82, n83, n84,
         n86, n88, n89, n90, n91, n92, n94, n96, n97, n98, n99, n100, n102,
         n104, n105, n106, n107, n108, n110, n112, n113, n114, n115, n116,
         n118, n120, n121, n122, n123, n124, n126, n128, n129, n130, n131,
         n133, n135, n136, n138, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n158,
         n160, n162, n164, n166, n168, n170, n172, n174, n176, n182, n184,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301;

  XOR2X1 U2 ( .A(B[31]), .B(A[31]), .Y(n1) );
  ADDFXL U3 ( .A(B[30]), .B(A[30]), .CI(n33), .CO(n32), .S(SUM[30]) );
  XOR2X1 U4 ( .A(n36), .B(n2), .Y(SUM[29]) );
  XOR2X1 U18 ( .A(n44), .B(n4), .Y(SUM[27]) );
  XOR2X1 U32 ( .A(n52), .B(n6), .Y(SUM[25]) );
  XOR2X1 U46 ( .A(n60), .B(n8), .Y(SUM[23]) );
  XOR2X1 U60 ( .A(n68), .B(n10), .Y(SUM[21]) );
  XOR2X1 U74 ( .A(n76), .B(n12), .Y(SUM[19]) );
  XOR2X1 U88 ( .A(n84), .B(n14), .Y(SUM[17]) );
  XOR2X1 U102 ( .A(n92), .B(n16), .Y(SUM[15]) );
  XOR2X1 U116 ( .A(n100), .B(n18), .Y(SUM[13]) );
  XOR2X1 U130 ( .A(n108), .B(n20), .Y(SUM[11]) );
  XOR2X1 U144 ( .A(n116), .B(n22), .Y(SUM[9]) );
  XOR2X1 U158 ( .A(n124), .B(n24), .Y(SUM[7]) );
  XOR2X1 U172 ( .A(n136), .B(n26), .Y(SUM[5]) );
  XOR2X1 U199 ( .A(n150), .B(n29), .Y(SUM[2]) );
  XOR2X1 U205 ( .A(n30), .B(n155), .Y(SUM[1]) );
  XNOR2XL U220 ( .A(n129), .B(n25), .Y(SUM[6]) );
  NOR2XL U221 ( .A(B[1]), .B(A[1]), .Y(n152) );
  OAI21XL U222 ( .A0(n36), .A1(n34), .B0(n35), .Y(n33) );
  NAND2BX1 U223 ( .AN(n148), .B(n149), .Y(n29) );
  AOI21XL U224 ( .A0(n141), .A1(n288), .B0(n138), .Y(n136) );
  NAND2BX1 U225 ( .AN(n122), .B(n123), .Y(n24) );
  XNOR2XL U226 ( .A(n121), .B(n23), .Y(SUM[8]) );
  AOI21XL U227 ( .A0(n129), .A1(n290), .B0(n126), .Y(n124) );
  AOI21XL U228 ( .A0(n121), .A1(n291), .B0(n118), .Y(n116) );
  AOI21XL U229 ( .A0(n113), .A1(n295), .B0(n110), .Y(n108) );
  AOI21XL U230 ( .A0(n105), .A1(n296), .B0(n102), .Y(n100) );
  AOI21XL U231 ( .A0(n97), .A1(n293), .B0(n94), .Y(n92) );
  AOI21XL U232 ( .A0(n89), .A1(n294), .B0(n86), .Y(n84) );
  AOI21XL U233 ( .A0(n81), .A1(n292), .B0(n78), .Y(n76) );
  AOI21XL U234 ( .A0(n73), .A1(n300), .B0(n70), .Y(n68) );
  AOI21XL U235 ( .A0(n65), .A1(n297), .B0(n62), .Y(n60) );
  AOI21XL U236 ( .A0(n57), .A1(n298), .B0(n54), .Y(n52) );
  AOI21XL U237 ( .A0(n49), .A1(n299), .B0(n46), .Y(n44) );
  AOI21XL U238 ( .A0(n151), .A1(n143), .B0(n144), .Y(n142) );
  XNOR2XL U239 ( .A(n41), .B(n3), .Y(SUM[28]) );
  XNOR2XL U240 ( .A(n65), .B(n9), .Y(SUM[22]) );
  XNOR2XL U241 ( .A(n57), .B(n7), .Y(SUM[24]) );
  XNOR2XL U242 ( .A(n49), .B(n5), .Y(SUM[26]) );
  XNOR2XL U243 ( .A(n81), .B(n13), .Y(SUM[18]) );
  XNOR2XL U244 ( .A(n97), .B(n17), .Y(SUM[14]) );
  XNOR2XL U245 ( .A(n89), .B(n15), .Y(SUM[16]) );
  XNOR2XL U246 ( .A(n73), .B(n11), .Y(SUM[20]) );
  XNOR2XL U247 ( .A(n113), .B(n21), .Y(SUM[10]) );
  XNOR2XL U248 ( .A(n105), .B(n19), .Y(SUM[12]) );
  INVXL U249 ( .A(n152), .Y(n184) );
  NOR2XL U250 ( .A(B[2]), .B(A[2]), .Y(n148) );
  NOR2XL U251 ( .A(B[3]), .B(A[3]), .Y(n145) );
  NAND2XL U252 ( .A(B[0]), .B(A[0]), .Y(n155) );
  OR2XL U253 ( .A(B[4]), .B(A[4]), .Y(n288) );
  OR2XL U254 ( .A(B[5]), .B(A[5]), .Y(n289) );
  NAND2XL U255 ( .A(B[2]), .B(A[2]), .Y(n149) );
  NAND2XL U256 ( .A(B[6]), .B(A[6]), .Y(n128) );
  NAND2XL U257 ( .A(B[5]), .B(A[5]), .Y(n135) );
  NAND2XL U258 ( .A(B[4]), .B(A[4]), .Y(n140) );
  NAND2XL U259 ( .A(B[3]), .B(A[3]), .Y(n146) );
  NAND2XL U260 ( .A(B[1]), .B(A[1]), .Y(n153) );
  OR2XL U261 ( .A(B[6]), .B(A[6]), .Y(n290) );
  XOR2XL U262 ( .A(n32), .B(n1), .Y(SUM[31]) );
  NAND2BXL U263 ( .AN(n154), .B(n155), .Y(n31) );
  NOR2XL U264 ( .A(B[0]), .B(A[0]), .Y(n154) );
  CLKINVX1 U265 ( .A(n142), .Y(n141) );
  CLKINVX1 U266 ( .A(n151), .Y(n150) );
  OAI21XL U267 ( .A0(n152), .A1(n155), .B0(n153), .Y(n151) );
  OAI21XL U268 ( .A0(n149), .A1(n145), .B0(n146), .Y(n144) );
  NOR2X1 U269 ( .A(n148), .B(n145), .Y(n143) );
  OAI21XL U270 ( .A0(n124), .A1(n122), .B0(n123), .Y(n121) );
  OAI21XL U271 ( .A0(n142), .A1(n130), .B0(n131), .Y(n129) );
  NAND2X1 U272 ( .A(n288), .B(n289), .Y(n130) );
  AOI21X1 U273 ( .A0(n289), .A1(n138), .B0(n133), .Y(n131) );
  CLKINVX1 U274 ( .A(n135), .Y(n133) );
  XNOR2X1 U275 ( .A(n141), .B(n27), .Y(SUM[4]) );
  NAND2X1 U276 ( .A(n288), .B(n140), .Y(n27) );
  NAND2X1 U277 ( .A(n290), .B(n128), .Y(n25) );
  NAND2X1 U278 ( .A(n291), .B(n120), .Y(n23) );
  CLKINVX1 U279 ( .A(n128), .Y(n126) );
  XNOR2X1 U280 ( .A(n147), .B(n28), .Y(SUM[3]) );
  NAND2X1 U281 ( .A(n182), .B(n146), .Y(n28) );
  OAI21XL U282 ( .A0(n150), .A1(n148), .B0(n149), .Y(n147) );
  CLKINVX1 U283 ( .A(n145), .Y(n182) );
  NAND2X1 U284 ( .A(n289), .B(n135), .Y(n26) );
  CLKINVX1 U285 ( .A(n140), .Y(n138) );
  NAND2X1 U286 ( .A(n156), .B(n35), .Y(n2) );
  OAI21XL U287 ( .A0(n84), .A1(n82), .B0(n83), .Y(n81) );
  OAI21XL U288 ( .A0(n52), .A1(n50), .B0(n51), .Y(n49) );
  OAI21XL U289 ( .A0(n116), .A1(n114), .B0(n115), .Y(n113) );
  OAI21XL U290 ( .A0(n76), .A1(n74), .B0(n75), .Y(n73) );
  OAI21XL U291 ( .A0(n44), .A1(n42), .B0(n43), .Y(n41) );
  OAI21XL U292 ( .A0(n108), .A1(n106), .B0(n107), .Y(n105) );
  OAI21XL U293 ( .A0(n100), .A1(n98), .B0(n99), .Y(n97) );
  OAI21XL U294 ( .A0(n68), .A1(n66), .B0(n67), .Y(n65) );
  OAI21XL U295 ( .A0(n92), .A1(n90), .B0(n91), .Y(n89) );
  OAI21XL U296 ( .A0(n60), .A1(n58), .B0(n59), .Y(n57) );
  CLKINVX1 U297 ( .A(n120), .Y(n118) );
  CLKINVX1 U298 ( .A(n112), .Y(n110) );
  CLKINVX1 U299 ( .A(n104), .Y(n102) );
  CLKINVX1 U300 ( .A(n96), .Y(n94) );
  CLKINVX1 U301 ( .A(n88), .Y(n86) );
  CLKINVX1 U302 ( .A(n80), .Y(n78) );
  CLKINVX1 U303 ( .A(n72), .Y(n70) );
  CLKINVX1 U304 ( .A(n64), .Y(n62) );
  CLKINVX1 U305 ( .A(n56), .Y(n54) );
  CLKINVX1 U306 ( .A(n48), .Y(n46) );
  AOI21X1 U307 ( .A0(n41), .A1(n301), .B0(n38), .Y(n36) );
  CLKINVX1 U308 ( .A(n40), .Y(n38) );
  NAND2X1 U309 ( .A(n170), .B(n91), .Y(n16) );
  NAND2X1 U310 ( .A(n168), .B(n83), .Y(n14) );
  NAND2X1 U311 ( .A(n166), .B(n75), .Y(n12) );
  NAND2X1 U312 ( .A(n164), .B(n67), .Y(n10) );
  NAND2X1 U313 ( .A(n162), .B(n59), .Y(n8) );
  NAND2X1 U314 ( .A(n160), .B(n51), .Y(n6) );
  NAND2X1 U315 ( .A(n158), .B(n43), .Y(n4) );
  NAND2X1 U316 ( .A(n300), .B(n72), .Y(n11) );
  NAND2X1 U317 ( .A(n301), .B(n40), .Y(n3) );
  NAND2X1 U318 ( .A(n294), .B(n88), .Y(n15) );
  NAND2X1 U319 ( .A(n292), .B(n80), .Y(n13) );
  NAND2X1 U320 ( .A(n297), .B(n64), .Y(n9) );
  NAND2X1 U321 ( .A(n298), .B(n56), .Y(n7) );
  NAND2X1 U322 ( .A(n299), .B(n48), .Y(n5) );
  NAND2X1 U323 ( .A(n176), .B(n115), .Y(n22) );
  NAND2X1 U324 ( .A(n174), .B(n107), .Y(n20) );
  NAND2X1 U325 ( .A(n172), .B(n99), .Y(n18) );
  CLKINVX1 U326 ( .A(n82), .Y(n168) );
  CLKINVX1 U327 ( .A(n50), .Y(n160) );
  CLKINVX1 U328 ( .A(n114), .Y(n176) );
  CLKINVX1 U329 ( .A(n74), .Y(n166) );
  CLKINVX1 U330 ( .A(n42), .Y(n158) );
  CLKINVX1 U331 ( .A(n106), .Y(n174) );
  CLKINVX1 U332 ( .A(n98), .Y(n172) );
  CLKINVX1 U333 ( .A(n66), .Y(n164) );
  CLKINVX1 U334 ( .A(n34), .Y(n156) );
  CLKINVX1 U335 ( .A(n90), .Y(n170) );
  CLKINVX1 U336 ( .A(n58), .Y(n162) );
  NAND2X1 U337 ( .A(n184), .B(n153), .Y(n30) );
  NAND2X1 U338 ( .A(n295), .B(n112), .Y(n21) );
  NAND2X1 U339 ( .A(n296), .B(n104), .Y(n19) );
  NAND2X1 U340 ( .A(n293), .B(n96), .Y(n17) );
  NOR2X1 U341 ( .A(B[7]), .B(A[7]), .Y(n122) );
  NAND2X1 U342 ( .A(B[7]), .B(A[7]), .Y(n123) );
  NAND2X1 U343 ( .A(B[8]), .B(A[8]), .Y(n120) );
  OR2X1 U344 ( .A(B[8]), .B(A[8]), .Y(n291) );
  NAND2X1 U345 ( .A(B[14]), .B(A[14]), .Y(n96) );
  NOR2X1 U346 ( .A(B[17]), .B(A[17]), .Y(n82) );
  NAND2X1 U347 ( .A(B[16]), .B(A[16]), .Y(n88) );
  NOR2X1 U348 ( .A(B[9]), .B(A[9]), .Y(n114) );
  NOR2X1 U349 ( .A(B[19]), .B(A[19]), .Y(n74) );
  NAND2X1 U350 ( .A(B[17]), .B(A[17]), .Y(n83) );
  NOR2X1 U351 ( .A(B[11]), .B(A[11]), .Y(n106) );
  NOR2X1 U352 ( .A(B[13]), .B(A[13]), .Y(n98) );
  NAND2X1 U353 ( .A(B[10]), .B(A[10]), .Y(n112) );
  NAND2X1 U354 ( .A(B[12]), .B(A[12]), .Y(n104) );
  NAND2X1 U355 ( .A(B[18]), .B(A[18]), .Y(n80) );
  NOR2X1 U356 ( .A(B[15]), .B(A[15]), .Y(n90) );
  NAND2X1 U357 ( .A(B[9]), .B(A[9]), .Y(n115) );
  NAND2X1 U358 ( .A(B[19]), .B(A[19]), .Y(n75) );
  NAND2X1 U359 ( .A(B[11]), .B(A[11]), .Y(n107) );
  NAND2X1 U360 ( .A(B[13]), .B(A[13]), .Y(n99) );
  NAND2X1 U361 ( .A(B[15]), .B(A[15]), .Y(n91) );
  OR2X1 U362 ( .A(B[18]), .B(A[18]), .Y(n292) );
  OR2X1 U363 ( .A(B[14]), .B(A[14]), .Y(n293) );
  OR2X1 U364 ( .A(B[16]), .B(A[16]), .Y(n294) );
  OR2X1 U365 ( .A(B[10]), .B(A[10]), .Y(n295) );
  OR2X1 U366 ( .A(B[12]), .B(A[12]), .Y(n296) );
  NAND2X1 U367 ( .A(B[22]), .B(A[22]), .Y(n64) );
  NOR2X1 U368 ( .A(B[25]), .B(A[25]), .Y(n50) );
  NAND2X1 U369 ( .A(B[24]), .B(A[24]), .Y(n56) );
  NOR2X1 U370 ( .A(B[27]), .B(A[27]), .Y(n42) );
  NAND2X1 U371 ( .A(B[25]), .B(A[25]), .Y(n51) );
  NOR2X1 U372 ( .A(B[21]), .B(A[21]), .Y(n66) );
  NOR2X1 U373 ( .A(B[29]), .B(A[29]), .Y(n34) );
  NAND2X1 U374 ( .A(B[26]), .B(A[26]), .Y(n48) );
  NAND2X1 U375 ( .A(B[20]), .B(A[20]), .Y(n72) );
  NAND2X1 U376 ( .A(B[28]), .B(A[28]), .Y(n40) );
  NOR2X1 U377 ( .A(B[23]), .B(A[23]), .Y(n58) );
  NAND2X1 U378 ( .A(B[27]), .B(A[27]), .Y(n43) );
  NAND2X1 U379 ( .A(B[21]), .B(A[21]), .Y(n67) );
  NAND2X1 U380 ( .A(B[29]), .B(A[29]), .Y(n35) );
  NAND2X1 U381 ( .A(B[23]), .B(A[23]), .Y(n59) );
  OR2X1 U382 ( .A(B[22]), .B(A[22]), .Y(n297) );
  OR2X1 U383 ( .A(B[24]), .B(A[24]), .Y(n298) );
  OR2X1 U384 ( .A(B[26]), .B(A[26]), .Y(n299) );
  OR2X1 U385 ( .A(B[20]), .B(A[20]), .Y(n300) );
  OR2X1 U386 ( .A(B[28]), .B(A[28]), .Y(n301) );
  CLKINVX1 U387 ( .A(n31), .Y(SUM[0]) );
endmodule


module ALU ( ALUin1_i, ALUin2_i, ALUctrl_i, ALUresult_o, ALUzero_o );
  input [31:0] ALUin1_i;
  input [31:0] ALUin2_i;
  input [2:0] ALUctrl_i;
  output [31:0] ALUresult_o;
  output ALUzero_o;
  wire   N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125,
         N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136,
         N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147,
         N148, N149, N150, N151, N152, N153, N154, N155, n147, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108;

  ALU_DW01_cmp6_0 r299 ( .A(ALUin1_i), .B(ALUin2_i), .TC(1'b1), .LT(N155), 
        .EQ(ALUzero_o) );
  ALU_DW01_sub_1 sub_411 ( .A(ALUin1_i), .B(ALUin2_i), .CI(1'b0), .DIFF({N154, 
        N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, 
        N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, 
        N129, N128, N127, N126, N125, N124, N123}) );
  ALU_DW01_add_1 add_410 ( .A(ALUin1_i), .B(ALUin2_i), .CI(1'b0), .SUM({N122, 
        N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, 
        N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, 
        N97, N96, N95, N94, N93, N92, N91}) );
  NOR3X2 U5 ( .A(ALUctrl_i[2]), .B(n28), .C(ALUctrl_i[0]), .Y(n1) );
  NOR3X1 U6 ( .A(n29), .B(n28), .C(ALUctrl_i[0]), .Y(n2) );
  NAND3X1 U7 ( .A(n22), .B(n23), .C(n24), .Y(ALUresult_o[8]) );
  AO22XL U8 ( .A0(N120), .A1(n1), .B0(N152), .B1(n2), .Y(n99) );
  NAND3XL U9 ( .A(ALUin2_i[5]), .B(n105), .C(ALUin1_i[5]), .Y(n4) );
  NAND3XL U10 ( .A(ALUin2_i[3]), .B(n105), .C(ALUin1_i[3]), .Y(n16) );
  NAND3XL U11 ( .A(ALUin2_i[4]), .B(n105), .C(ALUin1_i[4]), .Y(n7) );
  AO22XL U12 ( .A0(N121), .A1(n1), .B0(N153), .B1(n2), .Y(n102) );
  AO22XL U13 ( .A0(N119), .A1(n1), .B0(N151), .B1(n2), .Y(n96) );
  CLKINVX1 U14 ( .A(n31), .Y(n105) );
  NAND3XL U15 ( .A(ALUin2_i[6]), .B(ALUin1_i[6]), .C(n105), .Y(n25) );
  AO22XL U16 ( .A0(N122), .A1(n1), .B0(N154), .B1(n2), .Y(n106) );
  AOI32XL U17 ( .A0(ALUin2_i[0]), .A1(n105), .A2(ALUin1_i[0]), .B0(n3), .B1(
        n32), .Y(n33) );
  OR2XL U18 ( .A(ALUin2_i[0]), .B(ALUin1_i[0]), .Y(n32) );
  NOR2X1 U19 ( .A(n31), .B(n30), .Y(n3) );
  AND3XL U20 ( .A(ALUin2_i[1]), .B(n105), .C(ALUin1_i[1]), .Y(n38) );
  NAND3X1 U21 ( .A(n4), .B(n5), .C(n6), .Y(ALUresult_o[5]) );
  OAI21XL U22 ( .A0(ALUin2_i[5]), .A1(ALUin1_i[5]), .B0(n3), .Y(n5) );
  AOI22X1 U23 ( .A0(N96), .A1(n1), .B0(N128), .B1(n2), .Y(n6) );
  NAND3X1 U24 ( .A(n7), .B(n8), .C(n9), .Y(ALUresult_o[4]) );
  OAI21XL U25 ( .A0(ALUin2_i[4]), .A1(ALUin1_i[4]), .B0(n3), .Y(n8) );
  AOI22X1 U26 ( .A0(N95), .A1(n1), .B0(N127), .B1(n2), .Y(n9) );
  NAND3X1 U27 ( .A(n13), .B(n14), .C(n15), .Y(ALUresult_o[2]) );
  NAND3X1 U28 ( .A(ALUin2_i[2]), .B(n105), .C(ALUin1_i[2]), .Y(n13) );
  OAI21XL U29 ( .A0(ALUin2_i[2]), .A1(ALUin1_i[2]), .B0(n3), .Y(n14) );
  AOI22X1 U30 ( .A0(N93), .A1(n1), .B0(N125), .B1(n2), .Y(n15) );
  NAND3X1 U31 ( .A(n16), .B(n17), .C(n18), .Y(ALUresult_o[3]) );
  OAI21XL U32 ( .A0(ALUin2_i[3]), .A1(ALUin1_i[3]), .B0(n3), .Y(n17) );
  AOI22X1 U33 ( .A0(N94), .A1(n1), .B0(N126), .B1(n2), .Y(n18) );
  AO22X1 U34 ( .A0(N106), .A1(n1), .B0(N138), .B1(n2), .Y(n57) );
  AO22X1 U35 ( .A0(N108), .A1(n1), .B0(N140), .B1(n2), .Y(n63) );
  AO22X1 U36 ( .A0(N110), .A1(n1), .B0(N142), .B1(n2), .Y(n69) );
  AO22X1 U37 ( .A0(N112), .A1(n1), .B0(N144), .B1(n2), .Y(n75) );
  AO22X1 U38 ( .A0(N114), .A1(n1), .B0(N146), .B1(n2), .Y(n81) );
  AO22X1 U39 ( .A0(N116), .A1(n1), .B0(N148), .B1(n2), .Y(n87) );
  AO22X1 U40 ( .A0(N118), .A1(n1), .B0(N150), .B1(n2), .Y(n93) );
  AO22X1 U41 ( .A0(N111), .A1(n1), .B0(N143), .B1(n2), .Y(n72) );
  AO22X1 U42 ( .A0(N107), .A1(n1), .B0(N139), .B1(n2), .Y(n60) );
  AO22X1 U43 ( .A0(N109), .A1(n1), .B0(N141), .B1(n2), .Y(n66) );
  AO22X1 U44 ( .A0(N113), .A1(n1), .B0(N145), .B1(n2), .Y(n78) );
  AO22X1 U45 ( .A0(N115), .A1(n1), .B0(N147), .B1(n2), .Y(n84) );
  AO22X1 U46 ( .A0(N117), .A1(n1), .B0(N149), .B1(n2), .Y(n90) );
  AO22X1 U47 ( .A0(N100), .A1(n1), .B0(N132), .B1(n2), .Y(n39) );
  AO22X1 U48 ( .A0(N102), .A1(n1), .B0(N134), .B1(n2), .Y(n45) );
  AO22X1 U49 ( .A0(N104), .A1(n1), .B0(N136), .B1(n2), .Y(n51) );
  AO22X1 U50 ( .A0(N92), .A1(n1), .B0(N124), .B1(n2), .Y(n36) );
  AO22X1 U51 ( .A0(N101), .A1(n1), .B0(N133), .B1(n2), .Y(n42) );
  AO22X1 U52 ( .A0(N103), .A1(n1), .B0(N135), .B1(n2), .Y(n48) );
  AO22X1 U53 ( .A0(N105), .A1(n1), .B0(N137), .B1(n2), .Y(n54) );
  OA21XL U54 ( .A0(ALUin2_i[1]), .A1(ALUin1_i[1]), .B0(n3), .Y(n37) );
  OA21XL U55 ( .A0(ALUin2_i[30]), .A1(ALUin1_i[30]), .B0(n3), .Y(n103) );
  OA21XL U56 ( .A0(ALUin2_i[31]), .A1(ALUin1_i[31]), .B0(n3), .Y(n107) );
  OA21XL U57 ( .A0(ALUin2_i[18]), .A1(ALUin1_i[18]), .B0(n3), .Y(n67) );
  OA21XL U58 ( .A0(ALUin2_i[9]), .A1(ALUin1_i[9]), .B0(n3), .Y(n40) );
  OA21XL U59 ( .A0(ALUin2_i[10]), .A1(ALUin1_i[10]), .B0(n3), .Y(n43) );
  OA21XL U60 ( .A0(ALUin2_i[11]), .A1(ALUin1_i[11]), .B0(n3), .Y(n46) );
  OA21XL U61 ( .A0(ALUin2_i[12]), .A1(ALUin1_i[12]), .B0(n3), .Y(n49) );
  OA21XL U62 ( .A0(ALUin2_i[13]), .A1(ALUin1_i[13]), .B0(n3), .Y(n52) );
  OA21XL U63 ( .A0(ALUin2_i[19]), .A1(ALUin1_i[19]), .B0(n3), .Y(n70) );
  OA21XL U64 ( .A0(ALUin2_i[20]), .A1(ALUin1_i[20]), .B0(n3), .Y(n73) );
  OA21XL U65 ( .A0(ALUin2_i[21]), .A1(ALUin1_i[21]), .B0(n3), .Y(n76) );
  OA21XL U66 ( .A0(ALUin2_i[26]), .A1(ALUin1_i[26]), .B0(n3), .Y(n91) );
  OA21XL U67 ( .A0(ALUin2_i[27]), .A1(ALUin1_i[27]), .B0(n3), .Y(n94) );
  OA21XL U68 ( .A0(ALUin2_i[28]), .A1(ALUin1_i[28]), .B0(n3), .Y(n97) );
  OA21XL U69 ( .A0(ALUin2_i[29]), .A1(ALUin1_i[29]), .B0(n3), .Y(n100) );
  OA21XL U70 ( .A0(ALUin2_i[15]), .A1(ALUin1_i[15]), .B0(n3), .Y(n58) );
  OA21XL U71 ( .A0(ALUin2_i[23]), .A1(ALUin1_i[23]), .B0(n3), .Y(n82) );
  OA21XL U72 ( .A0(ALUin2_i[14]), .A1(ALUin1_i[14]), .B0(n3), .Y(n55) );
  OA21XL U73 ( .A0(ALUin2_i[16]), .A1(ALUin1_i[16]), .B0(n3), .Y(n61) );
  OA21XL U74 ( .A0(ALUin2_i[17]), .A1(ALUin1_i[17]), .B0(n3), .Y(n64) );
  OA21XL U75 ( .A0(ALUin2_i[22]), .A1(ALUin1_i[22]), .B0(n3), .Y(n79) );
  OA21XL U76 ( .A0(ALUin2_i[24]), .A1(ALUin1_i[24]), .B0(n3), .Y(n85) );
  OA21XL U77 ( .A0(ALUin2_i[25]), .A1(ALUin1_i[25]), .B0(n3), .Y(n88) );
  NAND3X1 U78 ( .A(n19), .B(n20), .C(n21), .Y(ALUresult_o[7]) );
  NAND3X1 U79 ( .A(ALUin2_i[7]), .B(ALUin1_i[7]), .C(n105), .Y(n19) );
  OAI21XL U80 ( .A0(ALUin2_i[7]), .A1(ALUin1_i[7]), .B0(n3), .Y(n20) );
  AOI22X1 U81 ( .A0(N98), .A1(n1), .B0(N130), .B1(n2), .Y(n21) );
  NAND3X1 U82 ( .A(ALUin2_i[8]), .B(ALUin1_i[8]), .C(n105), .Y(n22) );
  OAI21XL U83 ( .A0(ALUin2_i[8]), .A1(ALUin1_i[8]), .B0(n3), .Y(n23) );
  AOI22X1 U84 ( .A0(N99), .A1(n1), .B0(N131), .B1(n2), .Y(n24) );
  NAND3X1 U85 ( .A(n25), .B(n26), .C(n27), .Y(ALUresult_o[6]) );
  OAI21XL U86 ( .A0(ALUin2_i[6]), .A1(ALUin1_i[6]), .B0(n3), .Y(n26) );
  AOI22X1 U87 ( .A0(N97), .A1(n1), .B0(N129), .B1(n2), .Y(n27) );
  AND4X1 U88 ( .A(N155), .B(ALUctrl_i[2]), .C(ALUctrl_i[1]), .D(ALUctrl_i[0]), 
        .Y(n147) );
  OAI2BB1X1 U89 ( .A0N(N123), .A1N(n2), .B0(n33), .Y(n34) );
  OR2X1 U90 ( .A(ALUctrl_i[1]), .B(ALUctrl_i[2]), .Y(n31) );
  CLKINVX1 U91 ( .A(ALUctrl_i[2]), .Y(n29) );
  CLKINVX1 U92 ( .A(ALUctrl_i[0]), .Y(n30) );
  CLKINVX1 U93 ( .A(ALUctrl_i[1]), .Y(n28) );
  CLKINVX1 U94 ( .A(n35), .Y(ALUresult_o[0]) );
  AOI211X1 U95 ( .A0(N91), .A1(n1), .B0(n34), .C0(n147), .Y(n35) );
  OR3X2 U96 ( .A(n44), .B(n43), .C(n42), .Y(ALUresult_o[10]) );
  AND3X2 U97 ( .A(ALUin2_i[10]), .B(n105), .C(ALUin1_i[10]), .Y(n44) );
  OR3X2 U98 ( .A(n47), .B(n46), .C(n45), .Y(ALUresult_o[11]) );
  AND3X2 U99 ( .A(ALUin2_i[11]), .B(n105), .C(ALUin1_i[11]), .Y(n47) );
  OR3X2 U100 ( .A(n50), .B(n49), .C(n48), .Y(ALUresult_o[12]) );
  AND3X2 U101 ( .A(ALUin2_i[12]), .B(n105), .C(ALUin1_i[12]), .Y(n50) );
  OR3X2 U102 ( .A(n53), .B(n52), .C(n51), .Y(ALUresult_o[13]) );
  AND3X2 U103 ( .A(ALUin2_i[13]), .B(n105), .C(ALUin1_i[13]), .Y(n53) );
  OR3X2 U104 ( .A(n56), .B(n55), .C(n54), .Y(ALUresult_o[14]) );
  AND3X2 U105 ( .A(ALUin2_i[14]), .B(n105), .C(ALUin1_i[14]), .Y(n56) );
  OR3X2 U106 ( .A(n104), .B(n103), .C(n102), .Y(ALUresult_o[30]) );
  AND3X2 U107 ( .A(ALUin2_i[30]), .B(n105), .C(ALUin1_i[30]), .Y(n104) );
  OR3X2 U108 ( .A(n108), .B(n107), .C(n106), .Y(ALUresult_o[31]) );
  AND3X2 U109 ( .A(ALUin2_i[31]), .B(n105), .C(ALUin1_i[31]), .Y(n108) );
  OR3X2 U110 ( .A(n38), .B(n37), .C(n36), .Y(ALUresult_o[1]) );
  OR3X2 U111 ( .A(n59), .B(n58), .C(n57), .Y(ALUresult_o[15]) );
  AND3X2 U112 ( .A(ALUin2_i[15]), .B(n105), .C(ALUin1_i[15]), .Y(n59) );
  OR3X2 U113 ( .A(n62), .B(n61), .C(n60), .Y(ALUresult_o[16]) );
  AND3X2 U114 ( .A(ALUin2_i[16]), .B(n105), .C(ALUin1_i[16]), .Y(n62) );
  OR3X2 U115 ( .A(n65), .B(n64), .C(n63), .Y(ALUresult_o[17]) );
  AND3X2 U116 ( .A(ALUin2_i[17]), .B(n105), .C(ALUin1_i[17]), .Y(n65) );
  OR3X2 U117 ( .A(n68), .B(n67), .C(n66), .Y(ALUresult_o[18]) );
  AND3X2 U118 ( .A(ALUin2_i[18]), .B(n105), .C(ALUin1_i[18]), .Y(n68) );
  OR3X2 U119 ( .A(n71), .B(n70), .C(n69), .Y(ALUresult_o[19]) );
  AND3X2 U120 ( .A(ALUin2_i[19]), .B(n105), .C(ALUin1_i[19]), .Y(n71) );
  OR3X2 U121 ( .A(n74), .B(n73), .C(n72), .Y(ALUresult_o[20]) );
  AND3X2 U122 ( .A(ALUin2_i[20]), .B(n105), .C(ALUin1_i[20]), .Y(n74) );
  OR3X2 U123 ( .A(n77), .B(n76), .C(n75), .Y(ALUresult_o[21]) );
  AND3X2 U124 ( .A(ALUin2_i[21]), .B(n105), .C(ALUin1_i[21]), .Y(n77) );
  OR3X2 U125 ( .A(n80), .B(n79), .C(n78), .Y(ALUresult_o[22]) );
  AND3X2 U126 ( .A(ALUin2_i[22]), .B(n105), .C(ALUin1_i[22]), .Y(n80) );
  OR3X2 U127 ( .A(n83), .B(n82), .C(n81), .Y(ALUresult_o[23]) );
  AND3X2 U128 ( .A(ALUin2_i[23]), .B(n105), .C(ALUin1_i[23]), .Y(n83) );
  OR3X2 U129 ( .A(n86), .B(n85), .C(n84), .Y(ALUresult_o[24]) );
  AND3X2 U130 ( .A(ALUin2_i[24]), .B(n105), .C(ALUin1_i[24]), .Y(n86) );
  OR3X2 U131 ( .A(n89), .B(n88), .C(n87), .Y(ALUresult_o[25]) );
  AND3X2 U132 ( .A(ALUin2_i[25]), .B(n105), .C(ALUin1_i[25]), .Y(n89) );
  OR3X2 U133 ( .A(n92), .B(n91), .C(n90), .Y(ALUresult_o[26]) );
  AND3X2 U134 ( .A(ALUin2_i[26]), .B(n105), .C(ALUin1_i[26]), .Y(n92) );
  OR3X2 U135 ( .A(n95), .B(n94), .C(n93), .Y(ALUresult_o[27]) );
  AND3X2 U136 ( .A(ALUin2_i[27]), .B(n105), .C(ALUin1_i[27]), .Y(n95) );
  OR3X2 U137 ( .A(n98), .B(n97), .C(n96), .Y(ALUresult_o[28]) );
  AND3X2 U138 ( .A(ALUin2_i[28]), .B(n105), .C(ALUin1_i[28]), .Y(n98) );
  OR3X2 U139 ( .A(n101), .B(n100), .C(n99), .Y(ALUresult_o[29]) );
  AND3X2 U140 ( .A(ALUin2_i[29]), .B(n105), .C(ALUin1_i[29]), .Y(n101) );
  OR3X2 U141 ( .A(n41), .B(n40), .C(n39), .Y(ALUresult_o[9]) );
  AND3X2 U142 ( .A(ALUin2_i[9]), .B(n105), .C(ALUin1_i[9]), .Y(n41) );
endmodule


module Adder_0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [31:1] carry;

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  NAND2X2 U1 ( .A(A[30]), .B(carry[30]), .Y(n15) );
  XOR2XL U2 ( .A(n14), .B(carry[30]), .Y(SUM[30]) );
  AND2X2 U3 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XL U4 ( .A(n6), .B(carry[16]), .Y(SUM[16]) );
  XOR2X1 U5 ( .A(B[20]), .B(A[20]), .Y(n2) );
  XOR2X1 U6 ( .A(n2), .B(carry[20]), .Y(SUM[20]) );
  NAND2X1 U7 ( .A(A[20]), .B(carry[20]), .Y(n3) );
  NAND2X1 U8 ( .A(B[20]), .B(carry[20]), .Y(n4) );
  NAND2X1 U9 ( .A(B[20]), .B(A[20]), .Y(n5) );
  NAND3X1 U10 ( .A(n3), .B(n4), .C(n5), .Y(carry[21]) );
  XOR2X1 U11 ( .A(B[16]), .B(A[16]), .Y(n6) );
  NAND2X1 U12 ( .A(A[16]), .B(carry[16]), .Y(n7) );
  NAND2X1 U13 ( .A(B[16]), .B(carry[16]), .Y(n8) );
  NAND2X1 U14 ( .A(B[16]), .B(A[16]), .Y(n9) );
  NAND3X1 U15 ( .A(n7), .B(n8), .C(n9), .Y(carry[17]) );
  XOR2XL U16 ( .A(n10), .B(carry[28]), .Y(SUM[28]) );
  XOR2X1 U17 ( .A(B[28]), .B(A[28]), .Y(n10) );
  NAND2XL U18 ( .A(A[28]), .B(carry[28]), .Y(n11) );
  NAND2XL U19 ( .A(B[28]), .B(carry[28]), .Y(n12) );
  NAND2X1 U20 ( .A(B[28]), .B(A[28]), .Y(n13) );
  NAND3X1 U21 ( .A(n11), .B(n12), .C(n13), .Y(carry[29]) );
  XOR2X1 U22 ( .A(B[30]), .B(A[30]), .Y(n14) );
  NAND2XL U23 ( .A(B[30]), .B(carry[30]), .Y(n16) );
  NAND2X1 U24 ( .A(B[30]), .B(A[30]), .Y(n17) );
  NAND3X1 U25 ( .A(n15), .B(n16), .C(n17), .Y(carry[31]) );
  XOR2X1 U26 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Adder_0 ( data0_i, data1_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  output [31:0] data_o;


  Adder_0_DW01_add_0 add_454 ( .A(data0_i), .B(data1_i), .CI(1'b0), .SUM(
        data_o) );
endmodule


module Adder_1_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58;
  wire   [31:1] carry;

  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  XOR3X1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX4 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  NAND3X2 U1 ( .A(n27), .B(n28), .C(n29), .Y(carry[22]) );
  AND2X2 U2 ( .A(B[0]), .B(A[0]), .Y(n1) );
  NAND2X1 U3 ( .A(A[30]), .B(carry[30]), .Y(n3) );
  NAND2X1 U4 ( .A(B[30]), .B(carry[30]), .Y(n4) );
  NAND2X1 U5 ( .A(B[30]), .B(A[30]), .Y(n5) );
  NAND3X1 U6 ( .A(n3), .B(n4), .C(n5), .Y(carry[31]) );
  NAND3X1 U7 ( .A(n7), .B(n8), .C(n9), .Y(carry[12]) );
  XOR2XL U8 ( .A(B[30]), .B(A[30]), .Y(n2) );
  XOR2XL U9 ( .A(n2), .B(carry[30]), .Y(SUM[30]) );
  XOR2X1 U10 ( .A(B[11]), .B(A[11]), .Y(n6) );
  XOR2XL U11 ( .A(n6), .B(carry[11]), .Y(SUM[11]) );
  NAND2X1 U12 ( .A(A[11]), .B(carry[11]), .Y(n7) );
  NAND2X1 U13 ( .A(B[11]), .B(carry[11]), .Y(n8) );
  NAND2X1 U14 ( .A(B[11]), .B(A[11]), .Y(n9) );
  NAND2X1 U15 ( .A(B[19]), .B(carry[19]), .Y(n33) );
  INVXL U16 ( .A(A[28]), .Y(n35) );
  XOR2XL U17 ( .A(n10), .B(carry[12]), .Y(SUM[12]) );
  XOR2X1 U18 ( .A(B[12]), .B(A[12]), .Y(n10) );
  NAND2X1 U19 ( .A(A[12]), .B(carry[12]), .Y(n11) );
  NAND2X1 U20 ( .A(B[12]), .B(carry[12]), .Y(n12) );
  NAND2X1 U21 ( .A(B[12]), .B(A[12]), .Y(n13) );
  NAND3X1 U22 ( .A(n11), .B(n12), .C(n13), .Y(carry[13]) );
  XOR2XL U23 ( .A(B[4]), .B(carry[4]), .Y(n14) );
  XOR2X1 U24 ( .A(n14), .B(A[4]), .Y(SUM[4]) );
  NAND2X1 U25 ( .A(carry[4]), .B(A[4]), .Y(n15) );
  NAND2X1 U26 ( .A(B[4]), .B(A[4]), .Y(n16) );
  NAND2X1 U27 ( .A(B[4]), .B(carry[4]), .Y(n17) );
  NAND3X1 U28 ( .A(n15), .B(n16), .C(n17), .Y(carry[5]) );
  XOR2X1 U29 ( .A(B[15]), .B(A[15]), .Y(n18) );
  XOR2XL U30 ( .A(n18), .B(carry[15]), .Y(SUM[15]) );
  NAND2X1 U31 ( .A(A[15]), .B(carry[15]), .Y(n19) );
  NAND2X1 U32 ( .A(B[15]), .B(carry[15]), .Y(n20) );
  NAND2X1 U33 ( .A(B[15]), .B(A[15]), .Y(n21) );
  NAND3X1 U34 ( .A(n19), .B(n20), .C(n21), .Y(carry[16]) );
  INVX1 U35 ( .A(n46), .Y(n34) );
  XOR2XL U36 ( .A(B[28]), .B(carry[28]), .Y(n46) );
  XOR2XL U37 ( .A(B[21]), .B(A[21]), .Y(n26) );
  NAND2X1 U38 ( .A(A[21]), .B(carry[21]), .Y(n27) );
  NAND2X1 U39 ( .A(B[21]), .B(carry[21]), .Y(n28) );
  NAND2X1 U40 ( .A(B[21]), .B(A[21]), .Y(n29) );
  XOR2X1 U41 ( .A(B[2]), .B(A[2]), .Y(n22) );
  XOR2XL U42 ( .A(n22), .B(carry[2]), .Y(SUM[2]) );
  NAND2X1 U43 ( .A(A[2]), .B(carry[2]), .Y(n23) );
  NAND2X1 U44 ( .A(B[2]), .B(carry[2]), .Y(n24) );
  NAND2X1 U45 ( .A(B[2]), .B(A[2]), .Y(n25) );
  NAND3X1 U46 ( .A(n23), .B(n24), .C(n25), .Y(carry[3]) );
  XOR2XL U47 ( .A(n26), .B(carry[21]), .Y(SUM[21]) );
  XOR2XL U48 ( .A(B[19]), .B(carry[19]), .Y(n30) );
  XOR2X1 U49 ( .A(n30), .B(A[19]), .Y(SUM[19]) );
  NAND2X1 U50 ( .A(carry[19]), .B(A[19]), .Y(n31) );
  NAND2X1 U51 ( .A(B[19]), .B(A[19]), .Y(n32) );
  NAND3X1 U52 ( .A(n31), .B(n32), .C(n33), .Y(carry[20]) );
  NAND2XL U53 ( .A(n46), .B(n35), .Y(n36) );
  NAND2X1 U54 ( .A(n34), .B(A[28]), .Y(n37) );
  NAND2XL U55 ( .A(n36), .B(n37), .Y(SUM[28]) );
  XOR2X1 U56 ( .A(B[17]), .B(A[17]), .Y(n38) );
  XOR2XL U57 ( .A(n38), .B(carry[17]), .Y(SUM[17]) );
  NAND2X1 U58 ( .A(A[17]), .B(carry[17]), .Y(n39) );
  NAND2X1 U59 ( .A(B[17]), .B(carry[17]), .Y(n40) );
  NAND2X1 U60 ( .A(B[17]), .B(A[17]), .Y(n41) );
  NAND3X1 U61 ( .A(n39), .B(n40), .C(n41), .Y(carry[18]) );
  NAND2X1 U62 ( .A(carry[28]), .B(A[28]), .Y(n47) );
  NAND2X1 U63 ( .A(B[28]), .B(carry[28]), .Y(n49) );
  XOR2XL U64 ( .A(B[22]), .B(A[22]), .Y(n42) );
  XOR2XL U65 ( .A(n42), .B(carry[22]), .Y(SUM[22]) );
  NAND2X1 U66 ( .A(A[22]), .B(carry[22]), .Y(n43) );
  NAND2X1 U67 ( .A(B[22]), .B(carry[22]), .Y(n44) );
  NAND2X1 U68 ( .A(B[22]), .B(A[22]), .Y(n45) );
  NAND3X1 U69 ( .A(n43), .B(n44), .C(n45), .Y(carry[23]) );
  NAND2XL U70 ( .A(B[28]), .B(A[28]), .Y(n48) );
  NAND3X1 U71 ( .A(n47), .B(n48), .C(n49), .Y(carry[29]) );
  XOR2XL U72 ( .A(B[24]), .B(A[24]), .Y(n50) );
  XOR2XL U73 ( .A(n50), .B(carry[24]), .Y(SUM[24]) );
  NAND2X1 U74 ( .A(A[24]), .B(carry[24]), .Y(n51) );
  NAND2X1 U75 ( .A(B[24]), .B(carry[24]), .Y(n52) );
  NAND2X1 U76 ( .A(B[24]), .B(A[24]), .Y(n53) );
  NAND3X1 U77 ( .A(n51), .B(n52), .C(n53), .Y(carry[25]) );
  XOR2XL U78 ( .A(B[26]), .B(A[26]), .Y(n54) );
  XOR2XL U79 ( .A(n54), .B(carry[26]), .Y(SUM[26]) );
  NAND2X1 U80 ( .A(A[26]), .B(carry[26]), .Y(n55) );
  NAND2X1 U81 ( .A(B[26]), .B(carry[26]), .Y(n56) );
  NAND2X1 U82 ( .A(B[26]), .B(A[26]), .Y(n57) );
  NAND3X1 U83 ( .A(n55), .B(n56), .C(n57), .Y(carry[27]) );
  CLKINVX1 U84 ( .A(A[0]), .Y(n58) );
  XNOR2X1 U85 ( .A(B[0]), .B(n58), .Y(SUM[0]) );
endmodule


module Adder_1 ( data0_i, data1_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  output [31:0] data_o;


  Adder_1_DW01_add_0 add_454 ( .A(data0_i), .B(data1_i), .CI(1'b0), .SUM(
        data_o) );
endmodule


module MUX2_32b_5 ( data0_i, data1_i, sel_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  output [31:0] data_o;
  input sel_i;
  wire   n1, n2, n3, n4, n5, n6, n7;

  AO22X1 U1 ( .A0(data1_i[27]), .A1(sel_i), .B0(data0_i[27]), .B1(n5), .Y(
        data_o[27]) );
  AO22XL U2 ( .A0(data1_i[28]), .A1(sel_i), .B0(data0_i[28]), .B1(n5), .Y(
        data_o[28]) );
  AO22XL U3 ( .A0(data1_i[23]), .A1(sel_i), .B0(data0_i[23]), .B1(n5), .Y(
        data_o[23]) );
  CLKBUFX3 U4 ( .A(n7), .Y(n4) );
  CLKBUFX3 U5 ( .A(n7), .Y(n2) );
  CLKBUFX3 U6 ( .A(n7), .Y(n3) );
  CLKBUFX3 U7 ( .A(n7), .Y(n5) );
  CLKBUFX3 U8 ( .A(n7), .Y(n6) );
  CLKINVX1 U9 ( .A(n1), .Y(n7) );
  CLKBUFX3 U10 ( .A(sel_i), .Y(n1) );
  AO22X1 U11 ( .A0(data1_i[18]), .A1(sel_i), .B0(data0_i[18]), .B1(n5), .Y(
        data_o[18]) );
  AO22X1 U12 ( .A0(data1_i[19]), .A1(sel_i), .B0(data0_i[19]), .B1(n5), .Y(
        data_o[19]) );
  AO22X1 U13 ( .A0(data1_i[20]), .A1(n1), .B0(data0_i[20]), .B1(n5), .Y(
        data_o[20]) );
  AO22X1 U14 ( .A0(data1_i[21]), .A1(sel_i), .B0(data0_i[21]), .B1(n5), .Y(
        data_o[21]) );
  AO22X1 U15 ( .A0(data1_i[24]), .A1(sel_i), .B0(data0_i[24]), .B1(n5), .Y(
        data_o[24]) );
  AO22X1 U16 ( .A0(data1_i[26]), .A1(sel_i), .B0(data0_i[26]), .B1(n5), .Y(
        data_o[26]) );
  AO22X1 U17 ( .A0(data1_i[29]), .A1(sel_i), .B0(data0_i[29]), .B1(n5), .Y(
        data_o[29]) );
  AO22X1 U18 ( .A0(data1_i[31]), .A1(sel_i), .B0(data0_i[31]), .B1(n6), .Y(
        data_o[31]) );
  AO22X1 U19 ( .A0(data1_i[30]), .A1(sel_i), .B0(data0_i[30]), .B1(n6), .Y(
        data_o[30]) );
  AO22X1 U20 ( .A0(data1_i[14]), .A1(sel_i), .B0(data0_i[14]), .B1(n4), .Y(
        data_o[14]) );
  AO22X1 U21 ( .A0(data1_i[13]), .A1(sel_i), .B0(data0_i[13]), .B1(n4), .Y(
        data_o[13]) );
  AO22X1 U22 ( .A0(data1_i[4]), .A1(sel_i), .B0(data0_i[4]), .B1(n6), .Y(
        data_o[4]) );
  AO22X1 U23 ( .A0(data1_i[6]), .A1(sel_i), .B0(data0_i[6]), .B1(n6), .Y(
        data_o[6]) );
  AO22X1 U24 ( .A0(data1_i[7]), .A1(sel_i), .B0(data0_i[7]), .B1(n6), .Y(
        data_o[7]) );
  AO22X1 U25 ( .A0(data1_i[3]), .A1(sel_i), .B0(data0_i[3]), .B1(n6), .Y(
        data_o[3]) );
  AO22X1 U26 ( .A0(data1_i[11]), .A1(sel_i), .B0(data0_i[11]), .B1(n3), .Y(
        data_o[11]) );
  AO22X1 U27 ( .A0(data1_i[10]), .A1(sel_i), .B0(data0_i[10]), .B1(n2), .Y(
        data_o[10]) );
  AO22X1 U28 ( .A0(data1_i[12]), .A1(sel_i), .B0(data0_i[12]), .B1(n3), .Y(
        data_o[12]) );
  AO22X1 U29 ( .A0(data1_i[5]), .A1(sel_i), .B0(data0_i[5]), .B1(n6), .Y(
        data_o[5]) );
  AO22X1 U30 ( .A0(data1_i[8]), .A1(sel_i), .B0(data0_i[8]), .B1(n6), .Y(
        data_o[8]) );
  AO22X1 U31 ( .A0(data1_i[0]), .A1(sel_i), .B0(data0_i[0]), .B1(n2), .Y(
        data_o[0]) );
  AO22X1 U32 ( .A0(data1_i[1]), .A1(sel_i), .B0(data0_i[1]), .B1(n5), .Y(
        data_o[1]) );
  AO22X1 U33 ( .A0(data1_i[2]), .A1(sel_i), .B0(data0_i[2]), .B1(n5), .Y(
        data_o[2]) );
  AO22X1 U34 ( .A0(data1_i[15]), .A1(sel_i), .B0(data0_i[15]), .B1(n5), .Y(
        data_o[15]) );
  AO22X1 U35 ( .A0(data1_i[16]), .A1(sel_i), .B0(data0_i[16]), .B1(n5), .Y(
        data_o[16]) );
  AO22X1 U36 ( .A0(data1_i[17]), .A1(sel_i), .B0(data0_i[17]), .B1(n5), .Y(
        data_o[17]) );
  AO22X1 U37 ( .A0(data1_i[22]), .A1(sel_i), .B0(data0_i[22]), .B1(n5), .Y(
        data_o[22]) );
  AO22X1 U38 ( .A0(data1_i[25]), .A1(sel_i), .B0(data0_i[25]), .B1(n5), .Y(
        data_o[25]) );
  AO22X1 U39 ( .A0(sel_i), .A1(data1_i[9]), .B0(data0_i[9]), .B1(n6), .Y(
        data_o[9]) );
endmodule


module MUX2_32b_4 ( data0_i, data1_i, sel_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  output [31:0] data_o;
  input sel_i;
  wire   n1, n2, n3, n4, n5, n6, n7;

  AO22XL U1 ( .A0(data1_i[28]), .A1(sel_i), .B0(data0_i[28]), .B1(n5), .Y(
        data_o[28]) );
  AO22XL U2 ( .A0(data1_i[26]), .A1(n1), .B0(data0_i[26]), .B1(n5), .Y(
        data_o[26]) );
  AO22XL U3 ( .A0(data1_i[23]), .A1(sel_i), .B0(data0_i[23]), .B1(n5), .Y(
        data_o[23]) );
  AO22XL U4 ( .A0(data1_i[27]), .A1(n1), .B0(data0_i[27]), .B1(n5), .Y(
        data_o[27]) );
  AO22XL U5 ( .A0(data1_i[24]), .A1(sel_i), .B0(data0_i[24]), .B1(n5), .Y(
        data_o[24]) );
  AO22XL U6 ( .A0(data1_i[25]), .A1(n1), .B0(data0_i[25]), .B1(n5), .Y(
        data_o[25]) );
  AO22XL U7 ( .A0(data1_i[22]), .A1(sel_i), .B0(data0_i[22]), .B1(n5), .Y(
        data_o[22]) );
  CLKBUFX3 U8 ( .A(n7), .Y(n4) );
  CLKBUFX3 U9 ( .A(n4), .Y(n2) );
  CLKBUFX3 U10 ( .A(n7), .Y(n3) );
  CLKBUFX3 U11 ( .A(n7), .Y(n5) );
  CLKBUFX3 U12 ( .A(n7), .Y(n6) );
  AO22X1 U13 ( .A0(data1_i[18]), .A1(sel_i), .B0(data0_i[18]), .B1(n5), .Y(
        data_o[18]) );
  AO22X1 U14 ( .A0(data1_i[19]), .A1(n1), .B0(data0_i[19]), .B1(n5), .Y(
        data_o[19]) );
  AO22X1 U15 ( .A0(data1_i[20]), .A1(n1), .B0(data0_i[20]), .B1(n5), .Y(
        data_o[20]) );
  AO22X1 U16 ( .A0(data1_i[21]), .A1(sel_i), .B0(data0_i[21]), .B1(n5), .Y(
        data_o[21]) );
  AO22X1 U17 ( .A0(data1_i[29]), .A1(n1), .B0(data0_i[29]), .B1(n5), .Y(
        data_o[29]) );
  AO22X1 U18 ( .A0(data1_i[31]), .A1(n1), .B0(data0_i[31]), .B1(n6), .Y(
        data_o[31]) );
  AO22X1 U19 ( .A0(data1_i[30]), .A1(sel_i), .B0(data0_i[30]), .B1(n6), .Y(
        data_o[30]) );
  CLKINVX1 U20 ( .A(n1), .Y(n7) );
  AO22X1 U21 ( .A0(data1_i[14]), .A1(sel_i), .B0(data0_i[14]), .B1(n4), .Y(
        data_o[14]) );
  AO22X1 U22 ( .A0(data1_i[13]), .A1(n1), .B0(data0_i[13]), .B1(n4), .Y(
        data_o[13]) );
  AO22X1 U23 ( .A0(data1_i[4]), .A1(sel_i), .B0(data0_i[4]), .B1(n6), .Y(
        data_o[4]) );
  AO22X1 U24 ( .A0(data1_i[6]), .A1(n1), .B0(data0_i[6]), .B1(n6), .Y(
        data_o[6]) );
  AO22X1 U25 ( .A0(data1_i[7]), .A1(sel_i), .B0(data0_i[7]), .B1(n6), .Y(
        data_o[7]) );
  AO22X1 U26 ( .A0(data1_i[3]), .A1(n1), .B0(data0_i[3]), .B1(n6), .Y(
        data_o[3]) );
  AO22X1 U27 ( .A0(data1_i[11]), .A1(sel_i), .B0(data0_i[11]), .B1(n3), .Y(
        data_o[11]) );
  AO22X1 U28 ( .A0(data1_i[10]), .A1(n1), .B0(data0_i[10]), .B1(n2), .Y(
        data_o[10]) );
  AO22X1 U29 ( .A0(data1_i[12]), .A1(sel_i), .B0(data0_i[12]), .B1(n3), .Y(
        data_o[12]) );
  AO22X1 U30 ( .A0(data1_i[5]), .A1(sel_i), .B0(data0_i[5]), .B1(n6), .Y(
        data_o[5]) );
  AO22X1 U31 ( .A0(data1_i[8]), .A1(n1), .B0(data0_i[8]), .B1(n6), .Y(
        data_o[8]) );
  AO22X1 U32 ( .A0(data1_i[0]), .A1(n1), .B0(data0_i[0]), .B1(n2), .Y(
        data_o[0]) );
  AO22X1 U33 ( .A0(data1_i[1]), .A1(sel_i), .B0(data0_i[1]), .B1(n5), .Y(
        data_o[1]) );
  AO22X1 U34 ( .A0(data1_i[2]), .A1(n1), .B0(data0_i[2]), .B1(n5), .Y(
        data_o[2]) );
  AO22X1 U35 ( .A0(data1_i[15]), .A1(n1), .B0(data0_i[15]), .B1(n5), .Y(
        data_o[15]) );
  AO22X1 U36 ( .A0(data1_i[16]), .A1(sel_i), .B0(data0_i[16]), .B1(n5), .Y(
        data_o[16]) );
  AO22X1 U37 ( .A0(data1_i[17]), .A1(n1), .B0(data0_i[17]), .B1(n5), .Y(
        data_o[17]) );
  AO22X1 U38 ( .A0(sel_i), .A1(data1_i[9]), .B0(data0_i[9]), .B1(n6), .Y(
        data_o[9]) );
  CLKBUFX3 U39 ( .A(sel_i), .Y(n1) );
endmodule


module MUX2_32b_3 ( data0_i, data1_i, sel_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  output [31:0] data_o;
  input sel_i;
  wire   n1, n2, n3, n4, n5, n6, n7;

  AO22XL U1 ( .A0(data1_i[26]), .A1(sel_i), .B0(data0_i[26]), .B1(n5), .Y(
        data_o[26]) );
  AO22X1 U2 ( .A0(data1_i[23]), .A1(sel_i), .B0(data0_i[23]), .B1(n5), .Y(
        data_o[23]) );
  AO22XL U3 ( .A0(data1_i[27]), .A1(n1), .B0(data0_i[27]), .B1(n5), .Y(
        data_o[27]) );
  AO22XL U4 ( .A0(data1_i[24]), .A1(sel_i), .B0(data0_i[24]), .B1(n5), .Y(
        data_o[24]) );
  AO22XL U5 ( .A0(data1_i[25]), .A1(n1), .B0(data0_i[25]), .B1(n5), .Y(
        data_o[25]) );
  AO22XL U6 ( .A0(data1_i[22]), .A1(sel_i), .B0(data0_i[22]), .B1(n5), .Y(
        data_o[22]) );
  AO22XL U7 ( .A0(data1_i[1]), .A1(sel_i), .B0(data0_i[1]), .B1(n5), .Y(
        data_o[1]) );
  AO22XL U8 ( .A0(data1_i[2]), .A1(n1), .B0(data0_i[2]), .B1(n5), .Y(data_o[2]) );
  AO22XL U9 ( .A0(data1_i[0]), .A1(n1), .B0(data0_i[0]), .B1(n2), .Y(data_o[0]) );
  AO22XL U10 ( .A0(data1_i[3]), .A1(n1), .B0(data0_i[3]), .B1(n6), .Y(
        data_o[3]) );
  AO22XL U11 ( .A0(data1_i[4]), .A1(sel_i), .B0(data0_i[4]), .B1(n6), .Y(
        data_o[4]) );
  AO22XL U12 ( .A0(data1_i[5]), .A1(n1), .B0(data0_i[5]), .B1(n6), .Y(
        data_o[5]) );
  CLKBUFX3 U13 ( .A(n7), .Y(n4) );
  CLKBUFX3 U14 ( .A(n4), .Y(n2) );
  CLKBUFX3 U15 ( .A(n7), .Y(n3) );
  CLKBUFX3 U16 ( .A(n7), .Y(n5) );
  CLKBUFX3 U17 ( .A(n7), .Y(n6) );
  AO22X1 U18 ( .A0(data1_i[18]), .A1(sel_i), .B0(data0_i[18]), .B1(n5), .Y(
        data_o[18]) );
  AO22X1 U19 ( .A0(data1_i[19]), .A1(n1), .B0(data0_i[19]), .B1(n5), .Y(
        data_o[19]) );
  AO22X1 U20 ( .A0(data1_i[20]), .A1(n1), .B0(data0_i[20]), .B1(n5), .Y(
        data_o[20]) );
  AO22X1 U21 ( .A0(data1_i[21]), .A1(sel_i), .B0(data0_i[21]), .B1(n5), .Y(
        data_o[21]) );
  AO22X1 U22 ( .A0(data1_i[28]), .A1(n1), .B0(data0_i[28]), .B1(n5), .Y(
        data_o[28]) );
  AO22X1 U23 ( .A0(data1_i[29]), .A1(sel_i), .B0(data0_i[29]), .B1(n5), .Y(
        data_o[29]) );
  AO22X1 U24 ( .A0(data1_i[31]), .A1(sel_i), .B0(data0_i[31]), .B1(n6), .Y(
        data_o[31]) );
  AO22X1 U25 ( .A0(data1_i[30]), .A1(n1), .B0(data0_i[30]), .B1(n6), .Y(
        data_o[30]) );
  CLKINVX1 U26 ( .A(n1), .Y(n7) );
  AO22X1 U27 ( .A0(data1_i[14]), .A1(sel_i), .B0(data0_i[14]), .B1(n4), .Y(
        data_o[14]) );
  AO22X1 U28 ( .A0(data1_i[13]), .A1(n1), .B0(data0_i[13]), .B1(n4), .Y(
        data_o[13]) );
  AO22X1 U29 ( .A0(data1_i[6]), .A1(n1), .B0(data0_i[6]), .B1(n6), .Y(
        data_o[6]) );
  AO22X1 U30 ( .A0(data1_i[7]), .A1(sel_i), .B0(data0_i[7]), .B1(n6), .Y(
        data_o[7]) );
  AO22X1 U31 ( .A0(data1_i[11]), .A1(sel_i), .B0(data0_i[11]), .B1(n3), .Y(
        data_o[11]) );
  AO22X1 U32 ( .A0(data1_i[10]), .A1(n1), .B0(data0_i[10]), .B1(n2), .Y(
        data_o[10]) );
  AO22X1 U33 ( .A0(data1_i[12]), .A1(sel_i), .B0(data0_i[12]), .B1(n3), .Y(
        data_o[12]) );
  AO22X1 U34 ( .A0(data1_i[8]), .A1(n1), .B0(data0_i[8]), .B1(n6), .Y(
        data_o[8]) );
  AO22X1 U35 ( .A0(data1_i[15]), .A1(n1), .B0(data0_i[15]), .B1(n5), .Y(
        data_o[15]) );
  AO22X1 U36 ( .A0(data1_i[16]), .A1(sel_i), .B0(data0_i[16]), .B1(n5), .Y(
        data_o[16]) );
  AO22X1 U37 ( .A0(data1_i[17]), .A1(n1), .B0(data0_i[17]), .B1(n5), .Y(
        data_o[17]) );
  AO22X1 U38 ( .A0(sel_i), .A1(data1_i[9]), .B0(data0_i[9]), .B1(n6), .Y(
        data_o[9]) );
  CLKBUFX3 U39 ( .A(sel_i), .Y(n1) );
endmodule


module MUX2_32b_2 ( data0_i, data1_i, sel_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  output [31:0] data_o;
  input sel_i;
  wire   n1, n2, n3, n4, n5, n6, n7;

  AO22X1 U1 ( .A0(data1_i[28]), .A1(sel_i), .B0(data0_i[28]), .B1(n5), .Y(
        data_o[28]) );
  AO22X1 U2 ( .A0(data1_i[30]), .A1(n1), .B0(data0_i[30]), .B1(n6), .Y(
        data_o[30]) );
  AO22X1 U3 ( .A0(data1_i[29]), .A1(sel_i), .B0(data0_i[29]), .B1(n5), .Y(
        data_o[29]) );
  AO22X1 U4 ( .A0(data1_i[27]), .A1(n1), .B0(data0_i[27]), .B1(n5), .Y(
        data_o[27]) );
  AO22X1 U5 ( .A0(data1_i[31]), .A1(n1), .B0(data0_i[31]), .B1(n6), .Y(
        data_o[31]) );
  CLKBUFX3 U6 ( .A(n7), .Y(n4) );
  CLKBUFX3 U7 ( .A(n4), .Y(n2) );
  CLKBUFX3 U8 ( .A(n7), .Y(n3) );
  CLKBUFX3 U9 ( .A(n7), .Y(n5) );
  CLKBUFX3 U10 ( .A(n7), .Y(n6) );
  CLKINVX1 U11 ( .A(n1), .Y(n7) );
  CLKBUFX3 U12 ( .A(sel_i), .Y(n1) );
  AO22X1 U13 ( .A0(data1_i[0]), .A1(sel_i), .B0(data0_i[0]), .B1(n2), .Y(
        data_o[0]) );
  AO22X1 U14 ( .A0(data1_i[10]), .A1(n1), .B0(data0_i[10]), .B1(n2), .Y(
        data_o[10]) );
  AO22X1 U15 ( .A0(data1_i[11]), .A1(sel_i), .B0(data0_i[11]), .B1(n3), .Y(
        data_o[11]) );
  AO22X1 U16 ( .A0(data1_i[12]), .A1(n1), .B0(data0_i[12]), .B1(n3), .Y(
        data_o[12]) );
  AO22X1 U17 ( .A0(data1_i[13]), .A1(sel_i), .B0(data0_i[13]), .B1(n4), .Y(
        data_o[13]) );
  AO22X1 U18 ( .A0(data1_i[14]), .A1(n1), .B0(data0_i[14]), .B1(n4), .Y(
        data_o[14]) );
  AO22X1 U19 ( .A0(data1_i[3]), .A1(sel_i), .B0(data0_i[3]), .B1(n6), .Y(
        data_o[3]) );
  AO22X1 U20 ( .A0(data1_i[4]), .A1(n1), .B0(data0_i[4]), .B1(n6), .Y(
        data_o[4]) );
  AO22X1 U21 ( .A0(data1_i[5]), .A1(sel_i), .B0(data0_i[5]), .B1(n6), .Y(
        data_o[5]) );
  AO22X1 U22 ( .A0(data1_i[6]), .A1(n1), .B0(data0_i[6]), .B1(n6), .Y(
        data_o[6]) );
  AO22X1 U23 ( .A0(data1_i[7]), .A1(sel_i), .B0(data0_i[7]), .B1(n6), .Y(
        data_o[7]) );
  AO22X1 U24 ( .A0(data1_i[8]), .A1(n1), .B0(data0_i[8]), .B1(n6), .Y(
        data_o[8]) );
  AO22X1 U25 ( .A0(data1_i[1]), .A1(sel_i), .B0(data0_i[1]), .B1(n5), .Y(
        data_o[1]) );
  AO22X1 U26 ( .A0(data1_i[2]), .A1(sel_i), .B0(data0_i[2]), .B1(n5), .Y(
        data_o[2]) );
  AO22X1 U27 ( .A0(data1_i[15]), .A1(n1), .B0(data0_i[15]), .B1(n5), .Y(
        data_o[15]) );
  AO22X1 U28 ( .A0(data1_i[16]), .A1(sel_i), .B0(data0_i[16]), .B1(n5), .Y(
        data_o[16]) );
  AO22X1 U29 ( .A0(data1_i[17]), .A1(n1), .B0(data0_i[17]), .B1(n5), .Y(
        data_o[17]) );
  AO22X1 U30 ( .A0(data1_i[18]), .A1(sel_i), .B0(data0_i[18]), .B1(n5), .Y(
        data_o[18]) );
  AO22X1 U31 ( .A0(data1_i[19]), .A1(n1), .B0(data0_i[19]), .B1(n5), .Y(
        data_o[19]) );
  AO22X1 U32 ( .A0(data1_i[20]), .A1(n1), .B0(data0_i[20]), .B1(n5), .Y(
        data_o[20]) );
  AO22X1 U33 ( .A0(data1_i[21]), .A1(sel_i), .B0(data0_i[21]), .B1(n5), .Y(
        data_o[21]) );
  AO22X1 U34 ( .A0(data1_i[22]), .A1(n1), .B0(data0_i[22]), .B1(n5), .Y(
        data_o[22]) );
  AO22X1 U35 ( .A0(data1_i[23]), .A1(sel_i), .B0(data0_i[23]), .B1(n5), .Y(
        data_o[23]) );
  AO22X1 U36 ( .A0(data1_i[24]), .A1(n1), .B0(data0_i[24]), .B1(n5), .Y(
        data_o[24]) );
  AO22X1 U37 ( .A0(data1_i[25]), .A1(sel_i), .B0(data0_i[25]), .B1(n5), .Y(
        data_o[25]) );
  AO22X1 U38 ( .A0(data1_i[26]), .A1(n1), .B0(data0_i[26]), .B1(n5), .Y(
        data_o[26]) );
  AO22X1 U39 ( .A0(sel_i), .A1(data1_i[9]), .B0(data0_i[9]), .B1(n6), .Y(
        data_o[9]) );
endmodule


module MUX2_32b_1 ( data0_i, data1_i, sel_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  output [31:0] data_o;
  input sel_i;
  wire   n1, n2, n3, n4, n5, n6, n7;

  AO22XL U1 ( .A0(data1_i[28]), .A1(sel_i), .B0(data0_i[28]), .B1(n5), .Y(
        data_o[28]) );
  AO22XL U2 ( .A0(data1_i[29]), .A1(n1), .B0(data0_i[29]), .B1(n5), .Y(
        data_o[29]) );
  AO22XL U3 ( .A0(data1_i[30]), .A1(sel_i), .B0(data0_i[30]), .B1(n6), .Y(
        data_o[30]) );
  AO22X1 U4 ( .A0(data1_i[27]), .A1(sel_i), .B0(data0_i[27]), .B1(n5), .Y(
        data_o[27]) );
  AO22XL U5 ( .A0(data1_i[31]), .A1(n1), .B0(data0_i[31]), .B1(n6), .Y(
        data_o[31]) );
  AO22XL U6 ( .A0(data1_i[26]), .A1(n1), .B0(data0_i[26]), .B1(n5), .Y(
        data_o[26]) );
  AO22XL U7 ( .A0(data1_i[25]), .A1(sel_i), .B0(data0_i[25]), .B1(n5), .Y(
        data_o[25]) );
  AO22XL U8 ( .A0(data1_i[24]), .A1(n1), .B0(data0_i[24]), .B1(n5), .Y(
        data_o[24]) );
  AO22XL U9 ( .A0(data1_i[23]), .A1(sel_i), .B0(data0_i[23]), .B1(n5), .Y(
        data_o[23]) );
  AO22XL U10 ( .A0(data1_i[19]), .A1(n1), .B0(data0_i[19]), .B1(n5), .Y(
        data_o[19]) );
  AO22XL U11 ( .A0(data1_i[20]), .A1(n1), .B0(data0_i[20]), .B1(n5), .Y(
        data_o[20]) );
  AO22XL U12 ( .A0(data1_i[21]), .A1(sel_i), .B0(data0_i[21]), .B1(n5), .Y(
        data_o[21]) );
  AO22XL U13 ( .A0(data1_i[22]), .A1(n1), .B0(data0_i[22]), .B1(n5), .Y(
        data_o[22]) );
  AO22XL U14 ( .A0(data1_i[3]), .A1(n1), .B0(data0_i[3]), .B1(n6), .Y(
        data_o[3]) );
  AO22XL U15 ( .A0(data1_i[4]), .A1(n1), .B0(data0_i[4]), .B1(n6), .Y(
        data_o[4]) );
  AO22XL U16 ( .A0(data1_i[5]), .A1(n1), .B0(data0_i[5]), .B1(n6), .Y(
        data_o[5]) );
  AO22XL U17 ( .A0(data1_i[6]), .A1(n1), .B0(data0_i[6]), .B1(n6), .Y(
        data_o[6]) );
  AO22XL U18 ( .A0(data1_i[7]), .A1(n1), .B0(data0_i[7]), .B1(n6), .Y(
        data_o[7]) );
  AO22XL U19 ( .A0(data1_i[8]), .A1(sel_i), .B0(data0_i[8]), .B1(n6), .Y(
        data_o[8]) );
  AO22XL U20 ( .A0(data1_i[10]), .A1(sel_i), .B0(data0_i[10]), .B1(n2), .Y(
        data_o[10]) );
  AO22XL U21 ( .A0(data1_i[11]), .A1(n1), .B0(data0_i[11]), .B1(n3), .Y(
        data_o[11]) );
  AO22XL U22 ( .A0(data1_i[12]), .A1(sel_i), .B0(data0_i[12]), .B1(n3), .Y(
        data_o[12]) );
  AO22XL U23 ( .A0(data1_i[13]), .A1(n1), .B0(data0_i[13]), .B1(n4), .Y(
        data_o[13]) );
  AO22XL U24 ( .A0(data1_i[14]), .A1(sel_i), .B0(data0_i[14]), .B1(n4), .Y(
        data_o[14]) );
  AO22XL U25 ( .A0(data1_i[2]), .A1(sel_i), .B0(data0_i[2]), .B1(n5), .Y(
        data_o[2]) );
  AO22XL U26 ( .A0(data1_i[15]), .A1(n1), .B0(data0_i[15]), .B1(n5), .Y(
        data_o[15]) );
  AO22XL U27 ( .A0(data1_i[16]), .A1(n1), .B0(data0_i[16]), .B1(n5), .Y(
        data_o[16]) );
  AO22XL U28 ( .A0(data1_i[17]), .A1(sel_i), .B0(data0_i[17]), .B1(n5), .Y(
        data_o[17]) );
  AO22XL U29 ( .A0(data1_i[18]), .A1(n1), .B0(data0_i[18]), .B1(n5), .Y(
        data_o[18]) );
  CLKBUFX3 U30 ( .A(n7), .Y(n4) );
  CLKBUFX3 U31 ( .A(n4), .Y(n2) );
  CLKBUFX3 U32 ( .A(n7), .Y(n3) );
  CLKBUFX3 U33 ( .A(n7), .Y(n5) );
  CLKBUFX3 U34 ( .A(n7), .Y(n6) );
  CLKINVX1 U35 ( .A(n1), .Y(n7) );
  CLKBUFX3 U36 ( .A(sel_i), .Y(n1) );
  AO22X1 U37 ( .A0(data1_i[0]), .A1(n1), .B0(data0_i[0]), .B1(n2), .Y(
        data_o[0]) );
  AO22X1 U38 ( .A0(data1_i[1]), .A1(sel_i), .B0(data0_i[1]), .B1(n5), .Y(
        data_o[1]) );
  AO22X1 U39 ( .A0(n1), .A1(data1_i[9]), .B0(data0_i[9]), .B1(n6), .Y(
        data_o[9]) );
endmodule


module SingleCycle_MIPS ( clk, rst_n, IR_addr, IR, RF_writedata, ReadDataMem, 
        CEN, WEN, A, ReadData2, OEN );
  output [31:0] IR_addr;
  input [31:0] IR;
  output [31:0] RF_writedata;
  input [31:0] ReadDataMem;
  output [6:0] A;
  output [31:0] ReadData2;
  input clk, rst_n;
  output CEN, WEN, OEN;
  wire   RegDst, Jump, Branch, MemRead, MemToReg, MemWrite, ALUSrc, RegWrite,
         jal, jr, ALUresult_1, ALUresult_0, ALUzero, _3_net_, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17;
  wire   [31:0] PC_i;
  wire   [1:0] ALUOp;
  wire   [4:0] pre_Reg_W;
  wire   [4:0] Reg_W;
  wire   [31:0] ReadData1;
  wire   [31:0] IR_extend;
  wire   [31:0] ALUin2;
  wire   [2:0] ALUctrl;
  wire   [31:9] ALUresult;
  wire   [31:0] PC_add4;
  wire   [31:0] BranchAddr;
  wire   [31:0] MUX_Branch_o;
  wire   [31:0] MUX_Jump_o;
  wire   [31:0] MUX_MemToReg_o;
  assign OEN = 1'b0;

  PC PC ( .PC_i(PC_i), .PC_o(IR_addr), .clk(clk), .rst_n(n17) );
  Control Control ( .opcode_i(IR[31:26]), .func_i({IR[5:1], n6}), .RegDst_o(
        RegDst), .Jump_o(Jump), .Branch_o(Branch), .MemRead_o(MemRead), 
        .MemToReg_o(MemToReg), .ALUOp_o(ALUOp), .MemWrite_o(MemWrite), 
        .ALUSrc_o(ALUSrc), .RegWrite_o(RegWrite), .jal_o(jal), .jr_o(jr) );
  MUX2_5b_0 MUX_RegDST ( .data0_i({IR[20], n13, n12, n11, n10}), .data1_i(
        IR[15:11]), .sel_i(RegDst), .data_o(pre_Reg_W) );
  MUX2_5b_1 MUX_jal0 ( .data0_i(pre_Reg_W), .data1_i({1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1}), .sel_i(n8), .data_o(Reg_W) );
  Register Register ( .Reg_R1_i({IR[25], n16, IR[23], n15, n14}), .Reg_R2_i({
        IR[20], n13, n12, n11, n10}), .Reg_W_i(Reg_W), .RegWrite_i(RegWrite), 
        .WriteData_i(RF_writedata), .ReadData1_o(ReadData1), .ReadData2_o(
        ReadData2), .clk(clk), .rst_n(n17) );
  Sign_Extend Sign_Extend ( .data_i({IR[15:1], n6}), .data_o(IR_extend) );
  MUX2_32b_0 MUX_Src ( .data0_i(ReadData2), .data1_i(IR_extend), .sel_i(n9), 
        .data_o(ALUin2) );
  ALU_Control ALU_Control ( .func_i({IR[3:1], n7}), .ALUOp_i(ALUOp), 
        .ALUctrl_o(ALUctrl) );
  ALU ALU ( .ALUin1_i(ReadData1), .ALUin2_i(ALUin2), .ALUctrl_i(ALUctrl), 
        .ALUresult_o({ALUresult, A, ALUresult_1, ALUresult_0}), .ALUzero_o(
        ALUzero) );
  Adder_0 Adder0 ( .data0_i(IR_addr), .data1_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b0, 1'b0}), .data_o(PC_add4) );
  Adder_1 Adder1 ( .data0_i({PC_add4[31], n4, PC_add4[29:19], n3, 
        PC_add4[17:0]}), .data1_i({IR_extend[29:0], 1'b0, 1'b0}), .data_o(
        BranchAddr) );
  MUX2_32b_5 MUX_Branch ( .data0_i({PC_add4[31], n4, PC_add4[29:19], n3, 
        PC_add4[17:0]}), .data1_i(BranchAddr), .sel_i(_3_net_), .data_o(
        MUX_Branch_o) );
  MUX2_32b_4 MUX_Jump ( .data0_i(MUX_Branch_o), .data1_i({PC_add4[31], n4, 
        PC_add4[29:28], IR[25], n16, IR[23], n15, n14, IR[20], n13, n12, n11, 
        n10, IR[15:0], 1'b0, 1'b0}), .sel_i(Jump), .data_o(MUX_Jump_o) );
  MUX2_32b_3 MUX_jr ( .data0_i(MUX_Jump_o), .data1_i(ReadData1), .sel_i(jr), 
        .data_o(PC_i) );
  MUX2_32b_2 MUX_MemToReg ( .data0_i({ALUresult, A, ALUresult_1, ALUresult_0}), 
        .data1_i(ReadDataMem), .sel_i(MemToReg), .data_o(MUX_MemToReg_o) );
  MUX2_32b_1 MUX_jal1 ( .data0_i(MUX_MemToReg_o), .data1_i({PC_add4[31], n4, 
        PC_add4[29:19], n3, PC_add4[17:0]}), .sel_i(n8), .data_o(RF_writedata)
         );
  CLKINVX2 U7 ( .A(PC_add4[18]), .Y(n2) );
  INVX2 U8 ( .A(n2), .Y(n3) );
  BUFX3 U9 ( .A(PC_add4[30]), .Y(n4) );
  CLKINVX1 U10 ( .A(IR[0]), .Y(n5) );
  CLKINVX1 U11 ( .A(n5), .Y(n6) );
  CLKINVX1 U12 ( .A(n5), .Y(n7) );
  NOR2X1 U13 ( .A(MemWrite), .B(MemRead), .Y(CEN) );
  NAND2BX1 U14 ( .AN(MemRead), .B(MemWrite), .Y(WEN) );
  AND2X2 U15 ( .A(Branch), .B(ALUzero), .Y(_3_net_) );
  CLKBUFX3 U16 ( .A(jal), .Y(n8) );
  CLKBUFX3 U17 ( .A(ALUSrc), .Y(n9) );
  CLKBUFX3 U18 ( .A(rst_n), .Y(n17) );
  CLKBUFX3 U19 ( .A(IR[19]), .Y(n13) );
  CLKBUFX3 U20 ( .A(IR[18]), .Y(n12) );
  CLKBUFX3 U21 ( .A(IR[24]), .Y(n16) );
  CLKBUFX3 U22 ( .A(IR[16]), .Y(n10) );
  CLKBUFX3 U23 ( .A(IR[17]), .Y(n11) );
  CLKBUFX3 U24 ( .A(IR[21]), .Y(n14) );
  CLKBUFX3 U25 ( .A(IR[22]), .Y(n15) );
endmodule

